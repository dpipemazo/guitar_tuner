--
-- This is a test bench for the new sampling entity
--	Hopefully, maybe this thing will work.
--	That would be cool. I'm not terribly confident. 
--