/************************************************************************
 *                                                                      *
 * Copyright (c) 2009 Synfora, Inc.  All rights reserved.               *
 *                                                                      *
 * This file contains Confidential Information of Synfora, Inc.         *
 * In addition, certain inventions disclosed in this file may be        *
 * claimed within patents owned or patent applications filed by         *
 * Synfora or third parties.  Any use of Synfora's copyrighted works,   *
 * confidential information, patented inventions, or patent-pending     *
 * inventions is subject to the terms and conditions of your written    *
 * license agreement with Synfora, Inc.                                 *
 * All other use and disclosure is strictly prohibited.                 *
 *                                                                      *
 ************************************************************************/

/* Generated by PICO Extreme FPGA version 09.04 */
/* Target library : xilinx-spartan6-s2 */
/* Target frequency : 100 MHz */

`timescale 1ns / 10 ps
module test_pattern_generator_wide_ststream0_0_noreset(
        clk,
        reset,
        enable,
        flush,
        str_ready,
        sign,
        str_req,
        stallbar,
        pred,
        str_dataout,
        datain0,
        datain1,
        datain2,
        datain3,
        datain4,
        datain5);

  // Module parameters


  // synopsys template

  parameter sdwidth = 27;
  parameter strid = 0;
  parameter signwidth = 6;
  parameter dwidth0 = 8;
  parameter dwidth1 = 8;
  parameter dwidth2 = 8;
  parameter dwidth3 = 1;
  parameter dwidth4 = 1;
  parameter dwidth5 = 1;

  // Ports

  input  clk;
  input  reset;
  input  enable;
  input  flush;
  input  str_ready;
  input [signwidth - 1 : 0] sign;
  output  str_req;
  output  stallbar;
  input  pred;
  output [sdwidth - 1 : 0] str_dataout;
  input [dwidth0 - 1 : 0] datain0;
  input [dwidth1 - 1 : 0] datain1;
  input [dwidth2 - 1 : 0] datain2;
  input [dwidth3 - 1 : 0] datain3;
  input [dwidth4 - 1 : 0] datain4;
  input [dwidth5 - 1 : 0] datain5;

  // Wire/Reg for portformals 

  wire  clk;
  wire  reset;
  wire  enable;
  wire  flush;
  wire  str_ready;
  wire [signwidth - 1 : 0] sign;
  wire  str_req;
  wire  stallbar;
  wire  pred;
  wire [sdwidth - 1 : 0] str_dataout;
  wire [dwidth0 - 1 : 0] datain0;
  wire [dwidth1 - 1 : 0] datain1;
  wire [dwidth2 - 1 : 0] datain2;
  wire [dwidth3 - 1 : 0] datain3;
  wire [dwidth4 - 1 : 0] datain4;
  wire [dwidth5 - 1 : 0] datain5;


  // synopsys template

  parameter dwidth =   dwidth0+ dwidth1+ dwidth2+ dwidth3+ dwidth4+ dwidth5;

  parameter sdwidth0 = 8;

  parameter sdwidth1 = 8;

  parameter sdwidth2 = 8;

  parameter sdwidth3 = 1;

  parameter sdwidth4 = 1;

  parameter sdwidth5 = 1;

   // 0in assert -var (dwidth <= mdwidth)

  wire   [dwidth-1:0] st_packed_din;
  wire   [dwidth-1:0] st_packed_strout;

  wire   [sdwidth0+dwidth0-1:0] str_padded0;
  wire   [sdwidth1+dwidth1-1:0] str_padded1;
  wire   [sdwidth2+dwidth2-1:0] str_padded2;
  wire   [sdwidth3+dwidth3-1:0] str_padded3;
  wire   [sdwidth4+dwidth4-1:0] str_padded4;
  wire   [sdwidth5+dwidth5-1:0] str_padded5;

  assign st_packed_din[dwidth-1:0] = {
      datain5[dwidth5 - 1 : 0],
      datain4[dwidth4 - 1 : 0],
      datain3[dwidth3 - 1 : 0],
      datain2[dwidth2 - 1 : 0],
      datain1[dwidth1 - 1 : 0],
      datain0[dwidth0 - 1 : 0] };

	    assign str_padded0 = (sign[0]) ? {{sdwidth0{1'b0}}, st_packed_strout[0+dwidth0-1 : 0]} : {{sdwidth0{1'b0}} , st_packed_strout[0+dwidth0-1 : 0]};
  assign str_dataout[sdwidth0 + 0-1:0] = str_padded0[sdwidth0-1:0];
	    assign str_padded1 = (sign[1]) ? {{sdwidth1{1'b0}}, st_packed_strout[dwidth0 + 0+dwidth1-1 : dwidth0 + 0]} : {{sdwidth1{1'b0}} , st_packed_strout[dwidth0 + 0+dwidth1-1 : dwidth0 + 0]};
  assign str_dataout[sdwidth1 + sdwidth0 + 0-1:sdwidth0 + 0] = str_padded1[sdwidth1-1:0];
	    assign str_padded2 = (sign[2]) ? {{sdwidth2{1'b0}}, st_packed_strout[dwidth1 + dwidth0 + 0+dwidth2-1 : dwidth1 + dwidth0 + 0]} : {{sdwidth2{1'b0}} , st_packed_strout[dwidth1 + dwidth0 + 0+dwidth2-1 : dwidth1 + dwidth0 + 0]};
  assign str_dataout[sdwidth2 + sdwidth1 + sdwidth0 + 0-1:sdwidth1 + sdwidth0 + 0] = str_padded2[sdwidth2-1:0];
	    assign str_padded3 = (sign[3]) ? {{sdwidth3{1'b0}}, st_packed_strout[dwidth2 + dwidth1 + dwidth0 + 0+dwidth3-1 : dwidth2 + dwidth1 + dwidth0 + 0]} : {{sdwidth3{1'b0}} , st_packed_strout[dwidth2 + dwidth1 + dwidth0 + 0+dwidth3-1 : dwidth2 + dwidth1 + dwidth0 + 0]};
  assign str_dataout[sdwidth3 + sdwidth2 + sdwidth1 + sdwidth0 + 0-1:sdwidth2 + sdwidth1 + sdwidth0 + 0] = str_padded3[sdwidth3-1:0];
	    assign str_padded4 = (sign[4]) ? {{sdwidth4{1'b0}}, st_packed_strout[dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0+dwidth4-1 : dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0]} : {{sdwidth4{1'b0}} , st_packed_strout[dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0+dwidth4-1 : dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0]};
  assign str_dataout[sdwidth4 + sdwidth3 + sdwidth2 + sdwidth1 + sdwidth0 + 0-1:sdwidth3 + sdwidth2 + sdwidth1 + sdwidth0 + 0] = str_padded4[sdwidth4-1:0];
	    assign str_padded5 = (sign[5]) ? {{sdwidth5{1'b0}}, st_packed_strout[dwidth4 + dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0+dwidth5-1 : dwidth4 + dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0]} : {{sdwidth5{1'b0}} , st_packed_strout[dwidth4 + dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0+dwidth5-1 : dwidth4 + dwidth3 + dwidth2 + dwidth1 + dwidth0 + 0]};
  assign str_dataout[sdwidth5 + sdwidth4 + sdwidth3 + sdwidth2 + sdwidth1 + sdwidth0 + 0-1:sdwidth4 + sdwidth3 + sdwidth2 + sdwidth1 + sdwidth0 + 0] = str_padded5[sdwidth5-1:0];
  ststr_sx_noreset  #(.dwidth(dwidth), .sdwidth(dwidth), .strid(strid)) basic_instance(
      .enable(enable),
      .clk(clk),
      .reset(reset),
      .stallbar(stallbar),
      .flush(flush),
      .pred(pred),
      .str_req(str_req),
      .str_ready(str_ready),
      .sign(1'b0),
      .datain(st_packed_din),
      .str_dataout(st_packed_strout)
      );

endmodule


