/************************************************************************
 *                                                                      *
 * Copyright (c) 2009 Synfora, Inc.  All rights reserved.               *
 *                                                                      *
 * This file contains Confidential Information of Synfora, Inc.         *
 * In addition, certain inventions disclosed in this file may be        *
 * claimed within patents owned or patent applications filed by         *
 * Synfora or third parties.  Any use of Synfora's copyrighted works,   *
 * confidential information, patented inventions, or patent-pending     *
 * inventions is subject to the terms and conditions of your written    *
 * license agreement with Synfora, Inc.                                 *
 * All other use and disclosure is strictly prohibited.                 *
 *                                                                      *
 ************************************************************************/

/* Generated by PICO Extreme FPGA version 09.04 */
/* Target library : xilinx-spartan6-s2 */
/* Target frequency : 100 MHz */

`timescale 1ns / 10 ps
module test_pattern_generator(
        clk,
        reset,
        start_task_init,
        start_task_final,
        clear_init_done,
        clear_task_done,
        psw_livein_frames_in_use,
        psw_liveout_frames_in_use,
        psw_released,
        psw_sa_0_stalling,
        psw_busy,
        psw_idle,
        psw_init_done,
        psw_task_done,
        rawdatain_hsync_0,
        rawdatain_hblank_0,
        rawdatain_hbporch_0,
        rawdatain_hactive_0,
        rawdatain_vsync_0,
        rawdatain_vblank_0,
        rawdatain_vbporch_0,
        rawdatain_vactive_0,
        rawdatain_hfporch_0,
        rawdatain_vfporch_0,
        outstream_dvi_out_do_0_red,
        outstream_dvi_out_do_0_green,
        outstream_dvi_out_do_0_blue,
        outstream_dvi_out_do_0_hsync,
        outstream_dvi_out_do_0_vsync,
        outstream_dvi_out_do_0_de,
        outstream_dvi_out_req_0,
        outstream_dvi_out_ready_0);

  // Module parameters


  // synopsys template

  // Ports

  input  clk;
  input  reset;
  input  start_task_init;
  input  start_task_final;
  input  clear_init_done;
  input  clear_task_done;
  output [3 : 0] psw_livein_frames_in_use;
  output [3 : 0] psw_liveout_frames_in_use;
  output  psw_released;
  output  psw_sa_0_stalling;
  output  psw_busy;
  output  psw_idle;
  output  psw_init_done;
  output  psw_task_done;
  input  rawdatain_hsync_0;
  input [31 : 0] rawdatain_hblank_0;
  input [31 : 0] rawdatain_hbporch_0;
  input [31 : 0] rawdatain_hactive_0;
  input  rawdatain_vsync_0;
  input [31 : 0] rawdatain_vblank_0;
  input [31 : 0] rawdatain_vbporch_0;
  input [31 : 0] rawdatain_vactive_0;
  input [31 : 0] rawdatain_hfporch_0;
  input [31 : 0] rawdatain_vfporch_0;
  output [7 : 0] outstream_dvi_out_do_0_red;
  output [7 : 0] outstream_dvi_out_do_0_green;
  output [7 : 0] outstream_dvi_out_do_0_blue;
  output  outstream_dvi_out_do_0_hsync;
  output  outstream_dvi_out_do_0_vsync;
  output  outstream_dvi_out_do_0_de;
  output  outstream_dvi_out_req_0;
  input  outstream_dvi_out_ready_0;

  // Wire/Reg for portformals 

  wire  clk;
  wire  reset;
  wire  start_task_init;
  wire  start_task_final;
  wire  clear_init_done;
  wire  clear_task_done;
  wire [3 : 0] psw_livein_frames_in_use;
  wire [3 : 0] psw_liveout_frames_in_use;
  wire  psw_released;
  wire  psw_sa_0_stalling;
  wire  psw_busy;
  wire  psw_idle;
  wire  psw_init_done;
  wire  psw_task_done;
  wire  rawdatain_hsync_0;
  wire [31 : 0] rawdatain_hblank_0;
  wire [31 : 0] rawdatain_hbporch_0;
  wire [31 : 0] rawdatain_hactive_0;
  wire  rawdatain_vsync_0;
  wire [31 : 0] rawdatain_vblank_0;
  wire [31 : 0] rawdatain_vbporch_0;
  wire [31 : 0] rawdatain_vactive_0;
  wire [31 : 0] rawdatain_hfporch_0;
  wire [31 : 0] rawdatain_vfporch_0;
  wire [7 : 0] outstream_dvi_out_do_0_red;
  wire [7 : 0] outstream_dvi_out_do_0_green;
  wire [7 : 0] outstream_dvi_out_do_0_blue;
  wire  outstream_dvi_out_do_0_hsync;
  wire  outstream_dvi_out_do_0_vsync;
  wire  outstream_dvi_out_do_0_de;
  wire  outstream_dvi_out_req_0;
  wire  outstream_dvi_out_ready_0;

  wire [26 : 0] ppa_0_outstream_dvi_out_do_0;
  wire [26 : 0] combine8_wn_inst0_o0;
  wire [26 : 0] combine8_wn_inst1_o0;
  wire [26 : 0] combine8_wn_inst2_o0;


  // Signal assignments


  // Basic logic assignments


  // Component port and generic maps / Behavioural code.

  test_pattern_generator_ppa  ppa_0(
                      .clk(clk),
                      .reset(reset),
                      .start_task_init(start_task_init),
                      .start_task_final(start_task_final),
                      .clear_init_done(clear_init_done),
                      .clear_task_done(clear_task_done),
                      .psw_livein_frames_in_use(psw_livein_frames_in_use),
                      .psw_liveout_frames_in_use(psw_liveout_frames_in_use),
                      .psw_released(psw_released),
                      .psw_sa_0_stalling(psw_sa_0_stalling),
                      .psw_busy(psw_busy),
                      .psw_idle(psw_idle),
                      .psw_init_done(psw_init_done),
                      .psw_task_done(psw_task_done),
                      .rawdatain_hsync_0(rawdatain_hsync_0),
                      .rawdatain_hblank_0(rawdatain_hblank_0),
                      .rawdatain_hbporch_0(rawdatain_hbporch_0),
                      .rawdatain_hactive_0(rawdatain_hactive_0),
                      .rawdatain_vsync_0(rawdatain_vsync_0),
                      .rawdatain_vblank_0(rawdatain_vblank_0),
                      .rawdatain_vbporch_0(rawdatain_vbporch_0),
                      .rawdatain_vactive_0(rawdatain_vactive_0),
                      .rawdatain_hfporch_0(rawdatain_hfporch_0),
                      .rawdatain_vfporch_0(rawdatain_vfporch_0),
                      .outstream_dvi_out_do_0(ppa_0_outstream_dvi_out_do_0[26 : 0]),
                      .outstream_dvi_out_req_0(outstream_dvi_out_req_0),
                      .outstream_dvi_out_ready_0(outstream_dvi_out_ready_0));


  combine8_wn #(.inwidth(1))  combine8_wn_inst0(
                      .i0(ppa_0_outstream_dvi_out_do_0[0]),
                      .i1(ppa_0_outstream_dvi_out_do_0[1]),
                      .i2(ppa_0_outstream_dvi_out_do_0[2]),
                      .i3(ppa_0_outstream_dvi_out_do_0[3]),
                      .i4(ppa_0_outstream_dvi_out_do_0[4]),
                      .i5(ppa_0_outstream_dvi_out_do_0[5]),
                      .i6(ppa_0_outstream_dvi_out_do_0[6]),
                      .i7(ppa_0_outstream_dvi_out_do_0[7]),
                      .o0(combine8_wn_inst0_o0[7 : 0]));

  assign outstream_dvi_out_do_0_red = combine8_wn_inst0_o0[7 : 0];

  combine8_wn #(.inwidth(1))  combine8_wn_inst1(
                      .i0(ppa_0_outstream_dvi_out_do_0[8]),
                      .i1(ppa_0_outstream_dvi_out_do_0[9]),
                      .i2(ppa_0_outstream_dvi_out_do_0[10]),
                      .i3(ppa_0_outstream_dvi_out_do_0[11]),
                      .i4(ppa_0_outstream_dvi_out_do_0[12]),
                      .i5(ppa_0_outstream_dvi_out_do_0[13]),
                      .i6(ppa_0_outstream_dvi_out_do_0[14]),
                      .i7(ppa_0_outstream_dvi_out_do_0[15]),
                      .o0(combine8_wn_inst1_o0[7 : 0]));

  assign outstream_dvi_out_do_0_green = combine8_wn_inst1_o0[7 : 0];

  combine8_wn #(.inwidth(1))  combine8_wn_inst2(
                      .i0(ppa_0_outstream_dvi_out_do_0[16]),
                      .i1(ppa_0_outstream_dvi_out_do_0[17]),
                      .i2(ppa_0_outstream_dvi_out_do_0[18]),
                      .i3(ppa_0_outstream_dvi_out_do_0[19]),
                      .i4(ppa_0_outstream_dvi_out_do_0[20]),
                      .i5(ppa_0_outstream_dvi_out_do_0[21]),
                      .i6(ppa_0_outstream_dvi_out_do_0[22]),
                      .i7(ppa_0_outstream_dvi_out_do_0[23]),
                      .o0(combine8_wn_inst2_o0[7 : 0]));

  assign outstream_dvi_out_do_0_blue = combine8_wn_inst2_o0[7 : 0];
  assign outstream_dvi_out_do_0_hsync = ppa_0_outstream_dvi_out_do_0[24];
  assign outstream_dvi_out_do_0_vsync = ppa_0_outstream_dvi_out_do_0[25];
  assign outstream_dvi_out_do_0_de = ppa_0_outstream_dvi_out_do_0[26];


endmodule


