/************************************************************************
 *                                                                      *
 * Copyright (c) 2009 Synfora, Inc.  All rights reserved.               *
 *                                                                      *
 * This file contains Confidential Information of Synfora, Inc.         *
 * In addition, certain inventions disclosed in this file may be        *
 * claimed within patents owned or patent applications filed by         *
 * Synfora or third parties.  Any use of Synfora's copyrighted works,   *
 * confidential information, patented inventions, or patent-pending     *
 * inventions is subject to the terms and conditions of your written    *
 * license agreement with Synfora, Inc.                                 *
 * All other use and disclosure is strictly prohibited.                 *
 *                                                                      *
 ************************************************************************/

/* Generated by PICO Extreme FPGA version 09.04 */
/* Target library : xilinx-spartan6-s2 */
/* Target frequency : 100 MHz */

`timescale 1ns / 10 ps
module test_pattern_generator_pa_0(
        clk,
        reset,
        enable,
        start,
        abort,
        status,
        err,
        stallbar_in,
        stallbar_out,
        busy,
        outstream_dvi_out_do_0,
        outstream_dvi_out_req_0,
        outstream_dvi_out_ready_0,
        lid_rawdatain_hsync_0_0,
        lien_rawdatain_hsync_0_0,
        lid_rawdatain_hblank_0_0,
        lien_rawdatain_hblank_0_0,
        lid_rawdatain_hbporch_0_0,
        lien_rawdatain_hbporch_0_0,
        lid_rawdatain_hactive_0_0,
        lien_rawdatain_hactive_0_0,
        lid_rawdatain_vsync_0_0,
        lien_rawdatain_vsync_0_0,
        lid_rawdatain_vblank_0_0,
        lien_rawdatain_vblank_0_0,
        lid_rawdatain_vbporch_0_0,
        lien_rawdatain_vbporch_0_0,
        lid_rawdatain_vactive_0_0,
        lien_rawdatain_vactive_0_0,
        lid_rawdatain_hfporch_0_0,
        lien_rawdatain_hfporch_0_0,
        lid_rawdatain_vfporch_0_0,
        lien_rawdatain_vfporch_0_0);

  // Module parameters


  // synopsys template

  // Ports

  input  clk;
  input  reset;
  input  enable;
  input  start;
  input  abort;
  output  status;
  output  err;
  input  stallbar_in;
  output  stallbar_out;
  output  busy;
  output [26 : 0] outstream_dvi_out_do_0;
  output  outstream_dvi_out_req_0;
  input  outstream_dvi_out_ready_0;
  input  lid_rawdatain_hsync_0_0;
  input  lien_rawdatain_hsync_0_0;
  input [31 : 0] lid_rawdatain_hblank_0_0;
  input  lien_rawdatain_hblank_0_0;
  input [31 : 0] lid_rawdatain_hbporch_0_0;
  input  lien_rawdatain_hbporch_0_0;
  input [31 : 0] lid_rawdatain_hactive_0_0;
  input  lien_rawdatain_hactive_0_0;
  input  lid_rawdatain_vsync_0_0;
  input  lien_rawdatain_vsync_0_0;
  input [31 : 0] lid_rawdatain_vblank_0_0;
  input  lien_rawdatain_vblank_0_0;
  input [31 : 0] lid_rawdatain_vbporch_0_0;
  input  lien_rawdatain_vbporch_0_0;
  input [31 : 0] lid_rawdatain_vactive_0_0;
  input  lien_rawdatain_vactive_0_0;
  input [31 : 0] lid_rawdatain_hfporch_0_0;
  input  lien_rawdatain_hfporch_0_0;
  input [31 : 0] lid_rawdatain_vfporch_0_0;
  input  lien_rawdatain_vfporch_0_0;

  // Wire/Reg for portformals 

  wire  clk;
  wire  reset;
  wire  enable;
  wire  start;
  wire  abort;
  wire  status;
  wire  err;
  wire  stallbar_in;
  wire  stallbar_out;
  wire  busy;
  wire [26 : 0] outstream_dvi_out_do_0;
  wire  outstream_dvi_out_req_0;
  wire  outstream_dvi_out_ready_0;
  wire  lid_rawdatain_hsync_0_0;
  wire  lien_rawdatain_hsync_0_0;
  wire [31 : 0] lid_rawdatain_hblank_0_0;
  wire  lien_rawdatain_hblank_0_0;
  wire [31 : 0] lid_rawdatain_hbporch_0_0;
  wire  lien_rawdatain_hbporch_0_0;
  wire [31 : 0] lid_rawdatain_hactive_0_0;
  wire  lien_rawdatain_hactive_0_0;
  wire  lid_rawdatain_vsync_0_0;
  wire  lien_rawdatain_vsync_0_0;
  wire [31 : 0] lid_rawdatain_vblank_0_0;
  wire  lien_rawdatain_vblank_0_0;
  wire [31 : 0] lid_rawdatain_vbporch_0_0;
  wire  lien_rawdatain_vbporch_0_0;
  wire [31 : 0] lid_rawdatain_vactive_0_0;
  wire  lien_rawdatain_vactive_0_0;
  wire [31 : 0] lid_rawdatain_hfporch_0_0;
  wire  lien_rawdatain_hfporch_0_0;
  wire [31 : 0] lid_rawdatain_vfporch_0_0;
  wire  lien_rawdatain_vfporch_0_0;



  // Signal assignments


  // Basic logic assignments


  // Component port and generic maps / Behavioural code.

  test_pattern_generator_pe_0  pe_0(
                      .clk(clk),
                      .reset(reset),
                      .enable(enable),
                      .start(start),
                      .abort(abort),
                      .status(status),
                      .err(err),
                      .stallbar_in(stallbar_in),
                      .stallbar_out(stallbar_out),
                      .busy(busy),
                      .outstream_dvi_out_do_0(outstream_dvi_out_do_0),
                      .outstream_dvi_out_req_0(outstream_dvi_out_req_0),
                      .outstream_dvi_out_ready_0(outstream_dvi_out_ready_0),
                      .lid_rawdatain_hsync_0_0(lid_rawdatain_hsync_0_0),
                      .lien_rawdatain_hsync_0_0(lien_rawdatain_hsync_0_0),
                      .lid_rawdatain_hblank_0_0(lid_rawdatain_hblank_0_0),
                      .lien_rawdatain_hblank_0_0(lien_rawdatain_hblank_0_0),
                      .lid_rawdatain_hbporch_0_0(lid_rawdatain_hbporch_0_0),
                      .lien_rawdatain_hbporch_0_0(lien_rawdatain_hbporch_0_0),
                      .lid_rawdatain_hactive_0_0(lid_rawdatain_hactive_0_0),
                      .lien_rawdatain_hactive_0_0(lien_rawdatain_hactive_0_0),
                      .lid_rawdatain_vsync_0_0(lid_rawdatain_vsync_0_0),
                      .lien_rawdatain_vsync_0_0(lien_rawdatain_vsync_0_0),
                      .lid_rawdatain_vblank_0_0(lid_rawdatain_vblank_0_0),
                      .lien_rawdatain_vblank_0_0(lien_rawdatain_vblank_0_0),
                      .lid_rawdatain_vbporch_0_0(lid_rawdatain_vbporch_0_0),
                      .lien_rawdatain_vbporch_0_0(lien_rawdatain_vbporch_0_0),
                      .lid_rawdatain_vactive_0_0(lid_rawdatain_vactive_0_0),
                      .lien_rawdatain_vactive_0_0(lien_rawdatain_vactive_0_0),
                      .lid_rawdatain_hfporch_0_0(lid_rawdatain_hfporch_0_0),
                      .lien_rawdatain_hfporch_0_0(lien_rawdatain_hfporch_0_0),
                      .lid_rawdatain_vfporch_0_0(lid_rawdatain_vfporch_0_0),
                      .lien_rawdatain_vfporch_0_0(lien_rawdatain_vfporch_0_0));



endmodule


