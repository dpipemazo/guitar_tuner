/************************************************************************
 *                                                                      *
 * Copyright (c) 2009 Synfora, Inc.  All rights reserved.               *
 *                                                                      *
 * This file contains Confidential Information of Synfora, Inc.         *
 * In addition, certain inventions disclosed in this file may be        *
 * claimed within patents owned or patent applications filed by         *
 * Synfora or third parties.  Any use of Synfora's copyrighted works,   *
 * confidential information, patented inventions, or patent-pending     *
 * inventions is subject to the terms and conditions of your written    *
 * license agreement with Synfora, Inc.                                 *
 * All other use and disclosure is strictly prohibited.                 *
 *                                                                      *
 ************************************************************************/

/* Generated by PICO Extreme FPGA version 09.04 */
/* Target library : xilinx-spartan6-s2 */
/* Target frequency : 100 MHz */

`timescale 1ns / 10 ps
module test_pattern_generator_pe_0(
        clk,
        reset,
        enable,
        start,
        abort,
        status,
        err,
        stallbar_in,
        stallbar_out,
        busy,
        outstream_dvi_out_do_0,
        outstream_dvi_out_req_0,
        outstream_dvi_out_ready_0,
        lid_rawdatain_hsync_0_0,
        lien_rawdatain_hsync_0_0,
        lid_rawdatain_hblank_0_0,
        lien_rawdatain_hblank_0_0,
        lid_rawdatain_hbporch_0_0,
        lien_rawdatain_hbporch_0_0,
        lid_rawdatain_hactive_0_0,
        lien_rawdatain_hactive_0_0,
        lid_rawdatain_vsync_0_0,
        lien_rawdatain_vsync_0_0,
        lid_rawdatain_vblank_0_0,
        lien_rawdatain_vblank_0_0,
        lid_rawdatain_vbporch_0_0,
        lien_rawdatain_vbporch_0_0,
        lid_rawdatain_vactive_0_0,
        lien_rawdatain_vactive_0_0,
        lid_rawdatain_hfporch_0_0,
        lien_rawdatain_hfporch_0_0,
        lid_rawdatain_vfporch_0_0,
        lien_rawdatain_vfporch_0_0);

  // Module parameters


  // synopsys template

  // Ports

  input  clk;
  input  reset;
  input  enable;
  input  start;
  input  abort;
  output  status;
  output  err;
  input  stallbar_in;
  output  stallbar_out;
  output  busy;
  output [26 : 0] outstream_dvi_out_do_0;
  output  outstream_dvi_out_req_0;
  input  outstream_dvi_out_ready_0;
  input  lid_rawdatain_hsync_0_0;
  input  lien_rawdatain_hsync_0_0;
  input [31 : 0] lid_rawdatain_hblank_0_0;
  input  lien_rawdatain_hblank_0_0;
  input [31 : 0] lid_rawdatain_hbporch_0_0;
  input  lien_rawdatain_hbporch_0_0;
  input [31 : 0] lid_rawdatain_hactive_0_0;
  input  lien_rawdatain_hactive_0_0;
  input  lid_rawdatain_vsync_0_0;
  input  lien_rawdatain_vsync_0_0;
  input [31 : 0] lid_rawdatain_vblank_0_0;
  input  lien_rawdatain_vblank_0_0;
  input [31 : 0] lid_rawdatain_vbporch_0_0;
  input  lien_rawdatain_vbporch_0_0;
  input [31 : 0] lid_rawdatain_vactive_0_0;
  input  lien_rawdatain_vactive_0_0;
  input [31 : 0] lid_rawdatain_hfporch_0_0;
  input  lien_rawdatain_hfporch_0_0;
  input [31 : 0] lid_rawdatain_vfporch_0_0;
  input  lien_rawdatain_vfporch_0_0;

  // Wire/Reg for portformals 

  wire  clk;
  wire  reset;
  wire  enable;
  wire  start;
  wire  abort;
  wire  status;
  wire  err;
  wire  stallbar_in;
  wire  stallbar_out;
  wire  busy;
  wire [26 : 0] outstream_dvi_out_do_0;
  wire  outstream_dvi_out_req_0;
  wire  outstream_dvi_out_ready_0;
  wire  lid_rawdatain_hsync_0_0;
  wire  lien_rawdatain_hsync_0_0;
  wire [31 : 0] lid_rawdatain_hblank_0_0;
  wire  lien_rawdatain_hblank_0_0;
  wire [31 : 0] lid_rawdatain_hbporch_0_0;
  wire  lien_rawdatain_hbporch_0_0;
  wire [31 : 0] lid_rawdatain_hactive_0_0;
  wire  lien_rawdatain_hactive_0_0;
  wire  lid_rawdatain_vsync_0_0;
  wire  lien_rawdatain_vsync_0_0;
  wire [31 : 0] lid_rawdatain_vblank_0_0;
  wire  lien_rawdatain_vblank_0_0;
  wire [31 : 0] lid_rawdatain_vbporch_0_0;
  wire  lien_rawdatain_vbporch_0_0;
  wire [31 : 0] lid_rawdatain_vactive_0_0;
  wire  lien_rawdatain_vactive_0_0;
  wire [31 : 0] lid_rawdatain_hfporch_0_0;
  wire  lien_rawdatain_hfporch_0_0;
  wire [31 : 0] lid_rawdatain_vfporch_0_0;
  wire  lien_rawdatain_vfporch_0_0;

  wire  sig_enable;
  wire  sig_start;
  wire  sig_abort;
  wire  sig_stallbar_in;
  wire  inverter1n_inst42_o0;
  wire  or2n_inst2_o0;
  wire [26 : 0] outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_str_dataout;
  wire  outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_str_req;
  wire  sig_outstream_dvi_out_ready_0;
  wire  sig_lid_rawdatain_hsync_0_0;
  wire  sig_lien_rawdatain_hsync_0_0;
  wire [31 : 0] sig_lid_rawdatain_hblank_0_0;
  wire  sig_lien_rawdatain_hblank_0_0;
  wire [31 : 0] sig_lid_rawdatain_hbporch_0_0;
  wire  sig_lien_rawdatain_hbporch_0_0;
  wire [31 : 0] sig_lid_rawdatain_hactive_0_0;
  wire  sig_lien_rawdatain_hactive_0_0;
  wire  sig_lid_rawdatain_vsync_0_0;
  wire  sig_lien_rawdatain_vsync_0_0;
  wire [31 : 0] sig_lid_rawdatain_vblank_0_0;
  wire  sig_lien_rawdatain_vblank_0_0;
  wire [31 : 0] sig_lid_rawdatain_vbporch_0_0;
  wire  sig_lien_rawdatain_vbporch_0_0;
  wire [31 : 0] sig_lid_rawdatain_vactive_0_0;
  wire  sig_lien_rawdatain_vactive_0_0;
  wire [31 : 0] sig_lid_rawdatain_hfporch_0_0;
  wire  sig_lien_rawdatain_hfporch_0_0;
  wire [31 : 0] sig_lid_rawdatain_vfporch_0_0;
  wire  sig_lien_rawdatain_vfporch_0_0;
  wire  and3n_inst0_o0;
  wire  startbus;
  wire  and2n_inst0_o0;
  wire  and2n_inst2_o0;
  wire  controller_rsflipflop_noinit_inst0_q;
  wire  stagereg13_o0;
  wire  inverter1n_inst0_o0;
  wire  and2n_inst1_o0;
  wire  phasebus_0;
  wire  controller_rsflipflop_noinit_inst1_q;
  wire  or2n_inst1_o0;
  wire  and2n_inst8_o0;
  wire  and2n_inst3_o0;
  wire  and2n_inst4_o0;
  wire  and2n_inst6_o0;
  wire  and2n_inst5_o0;
  wire  inverter1n_inst1_o0;
  wire  and2n_inst7_o0;
  wire  stagereg1_o0;
  wire  stagereg2_o0;
  wire  stagereg3_o0;
  wire  stagereg4_o0;
  wire  stagereg5_o0;
  wire  stagereg6_o0;
  wire  stagereg7_o0;
  wire  stagereg8_o0;
  wire  stagereg9_o0;
  wire  stagereg10_o0;
  wire  stagereg11_o0;
  wire  stagereg12_o0;
  wire  delayed_done_o0;
  wire  rr_func_brf_inst0_stage_3_o0;
  wire [11 : 0] rr_var_x_stage_3_o0;
  wire [11 : 0] sext_inst16_o0;
  wire  cmpp_eq_inst0_o0_enable;
  wire  cmpp_eq_inst0_o0;
  wire  cmpp_eq_inst0_o1_enable;
  wire  cmpp_eq_inst0_o1;
  wire  rr_func_cmpp_eq_inst0_stage_6_o0;
  wire  sr_var_hsync_o0;
  wire  cmpp_eq_inst2_o0_enable;
  wire  cmpp_eq_inst2_o0;
  wire  cmpp_eq_inst2_o1_enable;
  wire  cmpp_eq_inst2_o1;
  wire  rr_func_cmpp_eq_inst0_0_stage_3_o0;
  wire [31 : 0] sext_inst4_o0;
  wire [31 : 0] sr_var_hblank_o0;
  wire  cmpp_eq_inst12_o0_enable;
  wire  cmpp_eq_inst12_o0;
  wire  cmpp_eq_inst12_o1_enable;
  wire  cmpp_eq_inst12_o1;
  wire  rr_func_cmpp_eq_inst12_stage_6_o0;
  wire  cmpp_eq_inst3_o0_enable;
  wire  cmpp_eq_inst3_o0;
  wire  cmpp_eq_inst3_o1_enable;
  wire  cmpp_eq_inst3_o1;
  wire  rr_func_cmpp_eq_inst12_0_stage_4_o0;
  wire [31 : 0] sr_var_hbporch_o0;
  wire  addw_inst4_o0_enable;
  wire [31 : 0] addw_inst4_o0;
  wire  rr_func_cmpp_eq_inst12_0_stage_5_o0;
  wire [31 : 0] sext_inst3_o0;
  wire [31 : 0] rr_func_addw_inst4_stage_5_o0;
  wire  cmpp_eq_inst13_o0_enable;
  wire  cmpp_eq_inst13_o0;
  wire  cmpp_eq_inst13_o1_enable;
  wire  cmpp_eq_inst13_o1;
  wire  rr_func_cmpp_eq_inst13_0_stage_6_o0;
  wire [31 : 0] rr_func_addw_inst4_stage_6_o0;
  wire [31 : 0] sr_var_hactive_1_o0;
  wire  addw_inst5_o0_enable;
  wire [31 : 0] addw_inst5_o0;
  wire  rr_func_cmpp_eq_inst13_0_stage_7_o0;
  wire [31 : 0] sext_inst2_o0;
  wire [31 : 0] rr_func_addw_inst5_stage_7_o0;
  wire  cmpp_eq_inst14_o0_enable;
  wire  cmpp_eq_inst14_o0;
  wire  cmpp_eq_inst14_o1_enable;
  wire  cmpp_eq_inst14_o1;
  wire  rr_func_brf_inst0_stage_7_o0;
  wire [11 : 0] rr_var_y_stage_7_o0;
  wire [11 : 0] sext_inst20_o0;
  wire  cmpp_eq_inst1_o0_enable;
  wire  cmpp_eq_inst1_o0;
  wire  cmpp_eq_inst1_o1_enable;
  wire  cmpp_eq_inst1_o1;
  wire  rr_func_cmpp_eq_inst1_stage_12_o0;
  wire  sr_var_vsync_o0;
  wire  cmpp_eq_inst4_o0_enable;
  wire  cmpp_eq_inst4_o0;
  wire  cmpp_eq_inst4_o1_enable;
  wire  cmpp_eq_inst4_o1;
  wire  rr_func_cmpp_eq_inst1_0_stage_7_o0;
  wire [31 : 0] sext_inst9_o0;
  wire [31 : 0] sr_var_vblank_o0;
  wire  cmpp_eq_inst15_o0_enable;
  wire  cmpp_eq_inst15_o0;
  wire  cmpp_eq_inst15_o1_enable;
  wire  cmpp_eq_inst15_o1;
  wire  rr_func_cmpp_eq_inst15_stage_12_o0;
  wire  cmpp_eq_inst5_o0_enable;
  wire  cmpp_eq_inst5_o0;
  wire  cmpp_eq_inst5_o1_enable;
  wire  cmpp_eq_inst5_o1;
  wire  rr_func_cmpp_eq_inst15_0_stage_8_o0;
  wire [31 : 0] sr_var_vbporch_o0;
  wire  addw_inst6_o0_enable;
  wire [31 : 0] addw_inst6_o0;
  wire  rr_func_cmpp_eq_inst15_0_stage_9_o0;
  wire [31 : 0] sext_inst8_o0;
  wire [31 : 0] rr_func_addw_inst6_stage_9_o0;
  wire  cmpp_eq_inst16_o0_enable;
  wire  cmpp_eq_inst16_o0;
  wire  cmpp_eq_inst16_o1_enable;
  wire  cmpp_eq_inst16_o1;
  wire  rr_func_cmpp_eq_inst16_0_stage_10_o0;
  wire [31 : 0] rr_func_addw_inst6_stage_10_o0;
  wire [31 : 0] sr_var_vactive_1_o0;
  wire  addw_inst7_o0_enable;
  wire [31 : 0] addw_inst7_o0;
  wire  rr_func_cmpp_eq_inst16_0_stage_11_o0;
  wire [31 : 0] sext_inst7_o0;
  wire [31 : 0] rr_func_addw_inst7_stage_11_o0;
  wire  cmpp_eq_inst17_o0_enable;
  wire  cmpp_eq_inst17_o0;
  wire  cmpp_eq_inst17_o1_enable;
  wire  cmpp_eq_inst17_o1;
  wire  rr_func_brf_inst0_stage_0_o0;
  wire  addw_inst8_o0_enable;
  wire [31 : 0] addw_inst8_o0;
  wire [31 : 0] sext_inst1_o0;
  wire [31 : 0] rr_func_addw_inst8_stage_2_o0;
  wire  cmpp_eq_inst18_o0_enable;
  wire  cmpp_eq_inst18_o0;
  wire  cmpp_eq_inst18_o1_enable;
  wire  cmpp_eq_inst18_o1;
  wire  rr_func_cmpp_eq_inst18_0_stage_3_o0;
  wire [32 : 0] sext_inst14_o0;
  wire  shrkw_inst0_o0_enable;
  wire [32 : 0] shrkw_inst0_o0;
  wire [28 : 0] sext_inst10_o0;
  wire  cmpp_eq_inst22_o0_enable;
  wire  cmpp_eq_inst22_o0;
  wire  cmpp_eq_inst22_o1_enable;
  wire  cmpp_eq_inst22_o1;
  wire  rr_func_cmpp_neq_inst0_0_stage_11_o0;
  wire [1 : 0] rr_var_ractive_stage_12_o0;
  wire [1 : 0] sext_inst27_o0;
  wire  cmpr_neq_inst1_o0_enable;
  wire [1 : 0] cmpr_neq_inst1_o0;
  wire [1 : 0] sext_inst28_o0;
  wire  cmpr_eq_inst1_o0_enable;
  wire [1 : 0] cmpr_eq_inst1_o0;
  wire  rr_func_cmpp_eq_inst22_stage_11_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst31_o0;
  wire [1 : 0] sext_inst29_o0;
  wire  cmpp_eq_inst6_o0_enable;
  wire  cmpp_eq_inst6_o0;
  wire  cmpp_eq_inst6_o1_enable;
  wire  cmpp_eq_inst6_o1;
  wire  rr_func_brf_inst0_stage_12_o0;
  wire [1 : 0] rr_var_gactive_stage_12_o0;
  wire [1 : 0] sext_inst30_o0;
  wire  cmpr_neq_inst2_o0_enable;
  wire [1 : 0] cmpr_neq_inst2_o0;
  wire [1 : 0] sext_inst31_o0;
  wire  cmpr_eq_inst2_o0_enable;
  wire [1 : 0] cmpr_eq_inst2_o0;
  wire [1 : 0] rr_var_bactive_stage_12_o0;
  wire [1 : 0] sext_inst32_o0;
  wire  cmpp_eq_inst7_o0_enable;
  wire  cmpp_eq_inst7_o0;
  wire  cmpp_eq_inst7_o1_enable;
  wire  cmpp_eq_inst7_o1;
  wire [1 : 0] sext_inst33_o0;
  wire  cmpr_neq_inst3_o0_enable;
  wire [1 : 0] cmpr_neq_inst3_o0;
  wire [1 : 0] sext_inst34_o0;
  wire  cmpr_eq_inst3_o0_enable;
  wire [1 : 0] cmpr_eq_inst3_o0;
  wire  rr_func_brf_inst0_stage_11_o0;
  wire [1 : 0] interconnect_select_3_1_wn_inst0_o0;
  wire [1 : 0] sext_inst35_o0;
  wire  cmpr_neq_inst0_o0_enable;
  wire [1 : 0] cmpr_neq_inst0_o0;
  wire [1 : 0] sext_inst36_o0;
  wire  cmpr_eq_inst0_o0_enable;
  wire [1 : 0] cmpr_eq_inst0_o0;
  wire  rr_func_cmpp_eq_inst22_stage_10_o0;
  wire [1 : 0] sext_inst37_o0;
  wire  cmpp_neq_inst0_o0_enable;
  wire  cmpp_neq_inst0_o0;
  wire  cmpp_neq_inst0_o1_enable;
  wire  cmpp_neq_inst0_o1;
  wire  rr_func_brf_inst0_stage_4_o0;
  wire [11 : 0] datamerge_select_2_1_wn_inst30_o0;
  wire [11 : 0] sext_inst38_o0;
  wire  addw_inst0_o0_enable;
  wire [11 : 0] addw_inst0_o0;
  wire  addw_inst9_o0_enable;
  wire [31 : 0] addw_inst9_o0;
  wire [31 : 0] sext_inst6_o0;
  wire [31 : 0] rr_func_addw_inst9_stage_6_o0;
  wire  cmpp_eq_inst19_o0_enable;
  wire  cmpp_eq_inst19_o0;
  wire  cmpp_eq_inst19_o1_enable;
  wire  cmpp_eq_inst19_o1;
  wire  rr_func_cmpp_eq_inst19_0_stage_7_o0;
  wire [32 : 0] sext_inst15_o0;
  wire  shrkw_inst1_o0_enable;
  wire [32 : 0] shrkw_inst1_o0;
  wire [30 : 0] sext_inst12_o0;
  wire  cmpp_eq_inst23_o0_enable;
  wire  cmpp_eq_inst23_o0;
  wire  cmpp_eq_inst23_o1_enable;
  wire  cmpp_eq_inst23_o1;
  wire  mpylw_multi_stage_noreset_inst0_o0_enable;
  wire [31 : 0] mpylw_multi_stage_noreset_inst0_o0;
  wire  rr_func_cmpp_eq_inst23_0_stage_8_o0;
  wire [32 : 0] sext_inst13_o0;
  wire  shrkw_inst2_o0_enable;
  wire [32 : 0] shrkw_inst2_o0;
  wire  rr_func_cmpp_eq_inst23_0_stage_9_o0;
  wire [29 : 0] sext_inst11_o0;
  wire [29 : 0] rr_func_shrkw_inst2_stage_9_o0;
  wire  cmpp_eq_inst24_o0_enable;
  wire  cmpp_eq_inst24_o0;
  wire  cmpp_eq_inst24_o1_enable;
  wire  cmpp_eq_inst24_o1;
  wire [1 : 0] datamerge_select_3_1_wn_inst8_o0;
  wire [1 : 0] sext_inst41_o0;
  wire  cmpp_neq_inst1_o0_enable;
  wire  cmpp_neq_inst1_o0;
  wire  cmpp_neq_inst1_o1_enable;
  wire  cmpp_neq_inst1_o1;
  wire  rr_func_cmpp_neq_inst1_stage_11_o0;
  wire [1 : 0] datamerge_select_3_1_wn_inst9_o0;
  wire [1 : 0] sext_inst42_o0;
  wire  cmpp_neq_inst2_o0_enable;
  wire  cmpp_neq_inst2_o0;
  wire  cmpp_neq_inst2_o1_enable;
  wire  cmpp_neq_inst2_o1;
  wire  rr_func_cmpp_neq_inst2_stage_12_o0;
  wire [1 : 0] sext_inst43_o0;
  wire  cmpr_neq_inst4_o0_enable;
  wire [1 : 0] cmpr_neq_inst4_o0;
  wire [1 : 0] datamerge_select_3_1_wn_inst5_o0;
  wire [1 : 0] sext_inst44_o0;
  wire  cmpp_eq_inst8_o0_enable;
  wire  cmpp_eq_inst8_o0;
  wire  cmpp_eq_inst8_o1_enable;
  wire  cmpp_eq_inst8_o1;
  wire [1 : 0] datamerge_select_3_1_wn_inst7_o0;
  wire [1 : 0] sext_inst45_o0;
  wire  cmpr_neq_inst5_o0_enable;
  wire [1 : 0] cmpr_neq_inst5_o0;
  wire  rr_func_cmpp_eq_inst8_0_stage_12_o0;
  wire [1 : 0] rr_func_cmpr_neq_inst5_stage_12_o0;
  wire [1 : 0] sext_inst46_o0;
  wire  cmpr_eq_inst4_o0_enable;
  wire [1 : 0] cmpr_eq_inst4_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst34_o0;
  wire [1 : 0] sext_inst47_o0;
  wire  cmpp_eq_inst9_o0_enable;
  wire  cmpp_eq_inst9_o0;
  wire  cmpp_eq_inst9_o1_enable;
  wire  cmpp_eq_inst9_o1;
  wire [1 : 0] datamerge_select_3_1_wn_inst6_o0;
  wire [1 : 0] sext_inst49_o0;
  wire  cmpr_neq_inst6_o0_enable;
  wire [1 : 0] cmpr_neq_inst6_o0;
  wire [1 : 0] rr_func_cmpr_neq_inst6_stage_12_o0;
  wire [1 : 0] sext_inst50_o0;
  wire  cmpr_eq_inst5_o0_enable;
  wire [1 : 0] cmpr_eq_inst5_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst36_o0;
  wire [1 : 0] sext_inst51_o0;
  wire  cmpp_eq_inst10_o0_enable;
  wire  cmpp_eq_inst10_o0;
  wire  cmpp_eq_inst10_o1_enable;
  wire  cmpp_eq_inst10_o1;
  wire  rr_func_cmpp_neq_inst2_0_stage_12_o0;
  wire [1 : 0] sext_inst53_o0;
  wire  cmpp_neq_inst3_o0_enable;
  wire  cmpp_neq_inst3_o0;
  wire  cmpp_neq_inst3_o1_enable;
  wire  cmpp_neq_inst3_o1;
  wire [1 : 0] sext_inst55_o0;
  wire  cmpp_neq_inst4_o0_enable;
  wire  cmpp_neq_inst4_o0;
  wire  cmpp_neq_inst4_o1_enable;
  wire  cmpp_neq_inst4_o1;
  wire  rr_func_cmpp_neq_inst1_stage_12_o0;
  wire [1 : 0] sext_inst57_o0;
  wire  cmpp_neq_inst5_o0_enable;
  wire  cmpp_neq_inst5_o0;
  wire  cmpp_neq_inst5_o1_enable;
  wire  cmpp_neq_inst5_o1;
  wire  rr_func_cmpp_neq_inst1_0_stage_12_o0;
  wire [1 : 0] sext_inst59_o0;
  wire  cmpp_neq_inst6_o0_enable;
  wire  cmpp_neq_inst6_o0;
  wire  cmpp_neq_inst6_o1_enable;
  wire  cmpp_neq_inst6_o1;
  wire  rr_func_brf_inst0_stage_13_o0;
  wire [1 : 0] datamerge_select_3_1_wn_inst2_o0;
  wire [1 : 0] sext_inst63_o0;
  wire  cmpr_neq_inst7_o0_enable;
  wire [1 : 0] cmpr_neq_inst7_o0;
  wire [1 : 0] sext_inst64_o0;
  wire  cmpp_eq_inst11_o0_enable;
  wire  cmpp_eq_inst11_o0;
  wire  cmpp_eq_inst11_o1_enable;
  wire  cmpp_eq_inst11_o1;
  wire [1 : 0] datamerge_select_3_1_wn_inst4_o0;
  wire [1 : 0] sext_inst65_o0;
  wire  cmpr_neq_inst8_o0_enable;
  wire [1 : 0] cmpr_neq_inst8_o0;
  wire  interconnect_select_1_1_wn_inst0_o0;
  wire [7 : 0] datamerge_select_3_1_wn_inst10_o0;
  wire [7 : 0] datamerge_select_3_1_wn_inst11_o0;
  wire [7 : 0] datamerge_select_2_1_wn_inst41_o0;
  wire  rr_var_dvi_ds_s_hs_stage_12_o0;
  wire  datamerge_select_3_1_wn_inst3_o0;
  wire [5 : 0] outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_combine6_wn_inst0_o0;
  wire  outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_stallbar;
  wire [31 : 0] sr_var_hfporch_o0;
  wire  addw_inst10_o0_enable;
  wire [31 : 0] addw_inst10_o0;
  wire  rr_func_brf_inst0_stage_1_o0;
  wire [31 : 0] rr_func_addw_inst8_stage_0_o0;
  wire [31 : 0] rr_func_addw_inst10_stage_0_o0;
  wire  addw_inst11_o0_enable;
  wire [31 : 0] addw_inst11_o0;
  wire  rr_func_brf_inst0_stage_2_o0;
  wire [31 : 0] rr_func_addw_inst11_stage_1_o0;
  wire [31 : 0] sext_inst66_o0;
  wire  addsubw_inst0_o0_enable;
  wire [31 : 0] addsubw_inst0_o0;
  wire [31 : 0] sext_inst0_o0;
  wire [31 : 0] rr_func_addsubw_inst0_stage_2_o0;
  wire  cmpp_eq_inst20_o0_enable;
  wire  cmpp_eq_inst20_o0;
  wire  cmpp_eq_inst20_o1_enable;
  wire  cmpp_eq_inst20_o1;
  wire  rr_func_cmpp_eq_inst20_stage_3_o0;
  wire [31 : 0] sr_var_vfporch_o0;
  wire  addw_inst12_o0_enable;
  wire [31 : 0] addw_inst12_o0;
  wire  rr_func_cmpp_eq_inst20_stage_4_o0;
  wire [31 : 0] rr_func_addw_inst9_stage_4_o0;
  wire [31 : 0] rr_func_addw_inst12_stage_4_o0;
  wire  addw_inst13_o0_enable;
  wire [31 : 0] addw_inst13_o0;
  wire  rr_func_cmpp_eq_inst20_stage_5_o0;
  wire [31 : 0] rr_func_addw_inst13_stage_5_o0;
  wire [31 : 0] sext_inst67_o0;
  wire  addsubw_inst1_o0_enable;
  wire [31 : 0] addsubw_inst1_o0;
  wire  rr_func_cmpp_eq_inst20_stage_6_o0;
  wire [31 : 0] sext_inst5_o0;
  wire [31 : 0] rr_func_addsubw_inst1_stage_6_o0;
  wire  cmpp_eq_inst21_o0_enable;
  wire  cmpp_eq_inst21_o0;
  wire  cmpp_eq_inst21_o1_enable;
  wire  cmpp_eq_inst21_o1;
  wire [11 : 0] sext_inst68_o0;
  wire  addw_inst1_o0_enable;
  wire [11 : 0] addw_inst1_o0;
  wire  rr_func_brf_inst0_stage_8_o0;
  wire [11 : 0] datamerge_select_2_1_wn_inst32_o0;
  wire [11 : 0] sext_inst69_o0;
  wire  addw_inst2_o0_enable;
  wire [11 : 0] addw_inst2_o0;
  wire [11 : 0] sext_inst70_o0;
  wire  addw_inst3_o0_enable;
  wire [11 : 0] addw_inst3_o0;
  wire  sr_var_loopcounter_o0;
  wire  brf_inst0_p_enable;
  wire  brf_inst0_p;
  wire  brf_inst0_lc_enable;
  wire  brf_inst0_lc_out;
  wire  brf_inst0_brf_o2_enable;
  wire  brf_inst0_brf_o2;
  wire  equal_inst0_o0;
  wire [11 : 0] rr_var_x_stage_8_o0;
  wire [11 : 0] rr_var_x_stage_6_o0;
  wire [11 : 0] rr_var_x_stage_4_o0;
  wire [11 : 0] rr_var_y_stage_12_o0;
  wire [11 : 0] rr_var_y_stage_10_o0;
  wire [11 : 0] rr_var_y_stage_8_o0;
  wire [1 : 0] sext_inst24_o0;
  wire  rr_func_cmpp_eq_inst18_stage_11_o0;
  wire  or2n_inst3_o0;
  wire [1 : 0] rr_func_moveii_inst40_stage_11_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_11_o0;
  wire  nor3n_inst0_o0;
  wire [11 : 0] rr_var_ya_1_stage_10_o0;
  wire [11 : 0] rr_var_ya_1_stage_8_o0;
  wire [1 : 0] sext_inst17_o0;
  wire [1 : 0] sext_inst18_o0;
  wire [1 : 0] sext_inst19_o0;
  wire [1 : 0] sext_inst21_o0;
  wire [1 : 0] sext_inst22_o0;
  wire [1 : 0] sext_inst23_o0;
  wire [1 : 0] sext_inst25_o0;
  wire [1 : 0] sext_inst26_o0;
  wire [1 : 0] sext_inst39_o0;
  wire [1 : 0] sext_inst40_o0;
  wire [8 : 0] sext_inst48_o0;
  wire [8 : 0] sext_inst52_o0;
  wire [8 : 0] sext_inst54_o0;
  wire [8 : 0] sext_inst56_o0;
  wire [8 : 0] sext_inst58_o0;
  wire [8 : 0] sext_inst60_o0;
  wire [8 : 0] sext_inst61_o0;
  wire [8 : 0] sext_inst62_o0;
  wire  and2n_inst9_o0;
  wire  or2n_inst4_o0;
  wire  select_2_1_wn_inst0_o0;
  wire  and2n_inst11_o0;
  wire  and2n_inst10_o0;
  wire  inverter1n_inst2_o0;
  wire  and2n_inst12_o0;
  wire  and2n_inst13_o0;
  wire  and2n_inst14_o0;
  wire  and2n_inst15_o0;
  wire  and2n_inst16_o0;
  wire  rr_func_brf_inst0_stage_5_o0;
  wire  and2n_inst17_o0;
  wire  rr_func_brf_inst0_stage_6_o0;
  wire  and2n_inst18_o0;
  wire  and2n_inst19_o0;
  wire  and2n_inst20_o0;
  wire  rr_func_brf_inst0_stage_9_o0;
  wire  and2n_inst21_o0;
  wire  rr_func_brf_inst0_stage_10_o0;
  wire  and2n_inst22_o0;
  wire  and2n_inst23_o0;
  wire  and2n_inst24_o0;
  wire  and2n_inst25_o0;
  wire  and2n_inst26_o0;
  wire  rr_func_cmpp_eq_inst0_stage_3_o0;
  wire  and2n_inst27_o0;
  wire  rr_func_cmpp_eq_inst0_stage_4_o0;
  wire  and2n_inst28_o0;
  wire  rr_func_cmpp_eq_inst0_stage_5_o0;
  wire  and2n_inst29_o0;
  wire  and2n_inst30_o0;
  wire  rr_func_cmpp_eq_inst0_stage_7_o0;
  wire  and2n_inst31_o0;
  wire  rr_func_cmpp_eq_inst0_stage_8_o0;
  wire  and2n_inst32_o0;
  wire  rr_func_cmpp_eq_inst0_stage_9_o0;
  wire  and2n_inst33_o0;
  wire  rr_func_cmpp_eq_inst0_stage_10_o0;
  wire  and2n_inst34_o0;
  wire  rr_func_cmpp_eq_inst0_stage_11_o0;
  wire  and2n_inst35_o0;
  wire  rr_func_cmpp_eq_inst0_stage_12_o0;
  wire  and2n_inst36_o0;
  wire  and2n_inst37_o0;
  wire  and2n_inst38_o0;
  wire  and2n_inst39_o0;
  wire  and2n_inst40_o0;
  wire  or3n_inst1_o0;
  wire  or2n_inst6_o0;
  wire  or3n_inst2_o0;
  wire  inverter1n_inst3_o0;
  wire [11 : 0] select_2_1_wn_inst1_o0;
  wire [11 : 0] select_2_1_wn_inst2_o0;
  wire  and2n_inst42_o0;
  wire [11 : 0] sext_inst71_o0;
  wire  and2n_inst44_o0;
  wire  and2n_inst41_o0;
  wire  inverter1n_inst4_o0;
  wire  or3n_inst3_o0;
  wire  and2n_inst43_o0;
  wire  inverter1n_inst5_o0;
  wire  and2n_inst45_o0;
  wire  and2n_inst46_o0;
  wire [11 : 0] rr_var_x_stage_5_o0;
  wire  and2n_inst47_o0;
  wire  and2n_inst48_o0;
  wire [11 : 0] rr_var_x_stage_7_o0;
  wire  and2n_inst49_o0;
  wire  and2n_inst50_o0;
  wire  and2n_inst51_o0;
  wire  or2n_inst9_o0;
  wire  or3n_inst4_o0;
  wire  inverter1n_inst6_o0;
  wire  select_2_1_wn_inst3_o0;
  wire  datamerge_select_2_1_wn_inst25_o0;
  wire  and2n_inst53_o0;
  wire  and2n_inst55_o0;
  wire  rr_var_dvi_ds_s_hs_stage_6_o0;
  wire  and2n_inst52_o0;
  wire  inverter1n_inst7_o0;
  wire  or2n_inst11_o0;
  wire  and3n_inst1_o0;
  wire  and2n_inst54_o0;
  wire  nor2n_inst0_o0;
  wire  nor2n_inst3_o0;
  wire  and2n_inst58_o0;
  wire  and2n_inst57_o0;
  wire  or2n_inst12_o0;
  wire  or2n_inst13_o0;
  wire  inverter1n_inst8_o0;
  wire  and2n_inst56_o0;
  wire  select_3_1_wn_inst1_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst26_o0;
  wire  and2n_inst59_o0;
  wire  rr_var_dvi_ds_s_hs_stage_7_o0;
  wire  and2n_inst60_o0;
  wire  rr_var_dvi_ds_s_hs_stage_8_o0;
  wire  and2n_inst61_o0;
  wire  rr_var_dvi_ds_s_hs_stage_9_o0;
  wire  and2n_inst62_o0;
  wire  rr_var_dvi_ds_s_hs_stage_10_o0;
  wire  and2n_inst63_o0;
  wire  rr_var_dvi_ds_s_hs_stage_11_o0;
  wire  and2n_inst64_o0;
  wire  and2n_inst65_o0;
  wire  and2n_inst66_o0;
  wire  rr_func_cmpp_eq_inst12_stage_4_o0;
  wire  and2n_inst67_o0;
  wire  rr_func_cmpp_eq_inst12_stage_5_o0;
  wire  and2n_inst68_o0;
  wire  and2n_inst69_o0;
  wire  rr_func_cmpp_eq_inst12_stage_7_o0;
  wire  and2n_inst70_o0;
  wire  rr_func_cmpp_eq_inst12_stage_8_o0;
  wire  and2n_inst71_o0;
  wire  rr_func_cmpp_eq_inst12_stage_9_o0;
  wire  and2n_inst72_o0;
  wire  rr_func_cmpp_eq_inst12_stage_10_o0;
  wire  and2n_inst73_o0;
  wire  rr_func_cmpp_eq_inst12_stage_11_o0;
  wire  and2n_inst74_o0;
  wire  rr_func_cmpp_eq_inst12_stage_12_o0;
  wire  and2n_inst75_o0;
  wire  and2n_inst76_o0;
  wire  and2n_inst77_o0;
  wire  and2n_inst78_o0;
  wire  and2n_inst79_o0;
  wire  and2n_inst80_o0;
  wire  and2n_inst81_o0;
  wire  and2n_inst82_o0;
  wire  rr_func_cmpp_eq_inst13_stage_6_o0;
  wire  and2n_inst83_o0;
  wire  rr_func_cmpp_eq_inst13_stage_7_o0;
  wire  and2n_inst84_o0;
  wire  rr_func_cmpp_eq_inst13_stage_8_o0;
  wire  and2n_inst85_o0;
  wire  rr_func_cmpp_eq_inst13_stage_9_o0;
  wire  and2n_inst86_o0;
  wire  rr_func_cmpp_eq_inst13_stage_10_o0;
  wire  and2n_inst87_o0;
  wire  rr_func_cmpp_eq_inst13_stage_11_o0;
  wire  and2n_inst88_o0;
  wire  rr_func_cmpp_eq_inst13_stage_12_o0;
  wire  and2n_inst89_o0;
  wire  and2n_inst90_o0;
  wire  and2n_inst91_o0;
  wire  or3n_inst6_o0;
  wire  or3n_inst7_o0;
  wire  and2n_inst92_o0;
  wire  and2n_inst93_o0;
  wire  and2n_inst94_o0;
  wire  and2n_inst95_o0;
  wire  and2n_inst96_o0;
  wire  and2n_inst97_o0;
  wire  or2n_inst14_o0;
  wire  or3n_inst8_o0;
  wire  or2n_inst15_o0;
  wire  or2n_inst16_o0;
  wire  or3n_inst9_o0;
  wire  inverter1n_inst9_o0;
  wire  rr_func_cmpp_eq_inst14_stage_12_o0;
  wire  rr_func_cmpp_eq_inst14_0_stage_12_o0;
  wire [1 : 0] select_2_1_wn_inst4_o0;
  wire [1 : 0] select_2_1_wn_inst5_o0;
  wire  and2n_inst99_o0;
  wire [1 : 0] sext_inst72_o0;
  wire  or3n_inst10_o0;
  wire  or2n_inst19_o0;
  wire  and2n_inst101_o0;
  wire [1 : 0] rr_var_hactive_stage_13_o0;
  wire  and2n_inst98_o0;
  wire  inverter1n_inst10_o0;
  wire  or3n_inst11_o0;
  wire  or3n_inst12_o0;
  wire  or2n_inst20_o0;
  wire  and2n_inst100_o0;
  wire  inverter1n_inst11_o0;
  wire  and2n_inst102_o0;
  wire  and2n_inst103_o0;
  wire  and2n_inst104_o0;
  wire  and2n_inst105_o0;
  wire  rr_func_cmpp_eq_inst14_stage_8_o0;
  wire  and2n_inst106_o0;
  wire  rr_func_cmpp_eq_inst14_stage_9_o0;
  wire  and2n_inst107_o0;
  wire  rr_func_cmpp_eq_inst14_stage_10_o0;
  wire  and2n_inst108_o0;
  wire  rr_func_cmpp_eq_inst14_stage_11_o0;
  wire  and2n_inst109_o0;
  wire  and2n_inst110_o0;
  wire  and2n_inst111_o0;
  wire  rr_func_cmpp_eq_inst14_0_stage_8_o0;
  wire  and2n_inst112_o0;
  wire  rr_func_cmpp_eq_inst14_0_stage_9_o0;
  wire  and2n_inst113_o0;
  wire  rr_func_cmpp_eq_inst14_0_stage_10_o0;
  wire  and2n_inst114_o0;
  wire  rr_func_cmpp_eq_inst14_0_stage_11_o0;
  wire  and2n_inst115_o0;
  wire  and2n_inst116_o0;
  wire  and2n_inst117_o0;
  wire  rr_func_cmpp_eq_inst1_stage_7_o0;
  wire  and2n_inst118_o0;
  wire  rr_func_cmpp_eq_inst1_stage_8_o0;
  wire  and2n_inst119_o0;
  wire  rr_func_cmpp_eq_inst1_stage_9_o0;
  wire  and2n_inst120_o0;
  wire  rr_func_cmpp_eq_inst1_stage_10_o0;
  wire  and2n_inst121_o0;
  wire  rr_func_cmpp_eq_inst1_stage_11_o0;
  wire  and2n_inst122_o0;
  wire  and2n_inst123_o0;
  wire  and2n_inst124_o0;
  wire  or3n_inst13_o0;
  wire  and2n_inst125_o0;
  wire  and2n_inst126_o0;
  wire  and2n_inst127_o0;
  wire  and2n_inst128_o0;
  wire  or2n_inst21_o0;
  wire  or3n_inst14_o0;
  wire  or3n_inst15_o0;
  wire  inverter1n_inst12_o0;
  wire  rr_func_cmpp_eq_inst20_0_stage_6_o0;
  wire [11 : 0] select_2_1_wn_inst6_o0;
  wire [11 : 0] select_2_1_wn_inst7_o0;
  wire  and2n_inst130_o0;
  wire [11 : 0] sext_inst73_o0;
  wire  or2n_inst24_o0;
  wire  and2n_inst132_o0;
  wire  and2n_inst129_o0;
  wire  inverter1n_inst13_o0;
  wire  or3n_inst16_o0;
  wire  or2n_inst25_o0;
  wire  and2n_inst131_o0;
  wire  inverter1n_inst14_o0;
  wire  and2n_inst133_o0;
  wire  and2n_inst134_o0;
  wire [11 : 0] rr_var_y_stage_9_o0;
  wire  and2n_inst135_o0;
  wire  and2n_inst136_o0;
  wire [11 : 0] rr_var_y_stage_11_o0;
  wire  and2n_inst137_o0;
  wire  and2n_inst138_o0;
  wire  and2n_inst139_o0;
  wire  or2n_inst26_o0;
  wire  or3n_inst17_o0;
  wire  inverter1n_inst15_o0;
  wire  rr_func_cmpp_eq_inst15_0_stage_11_o0;
  wire  select_2_1_wn_inst8_o0;
  wire  datamerge_select_2_1_wn_inst28_o0;
  wire  and2n_inst141_o0;
  wire  and2n_inst143_o0;
  wire  rr_var_dvi_ds_s_vs_stage_12_o0;
  wire  and2n_inst140_o0;
  wire  inverter1n_inst16_o0;
  wire  or2n_inst28_o0;
  wire  and3n_inst2_o0;
  wire  and2n_inst142_o0;
  wire  nor2n_inst1_o0;
  wire  nor2n_inst5_o0;
  wire  and2n_inst144_o0;
  wire  and2n_inst145_o0;
  wire  rr_func_cmpp_eq_inst15_stage_8_o0;
  wire  and2n_inst146_o0;
  wire  rr_func_cmpp_eq_inst15_stage_9_o0;
  wire  and2n_inst147_o0;
  wire  rr_func_cmpp_eq_inst15_stage_10_o0;
  wire  and2n_inst148_o0;
  wire  rr_func_cmpp_eq_inst15_stage_11_o0;
  wire  and2n_inst149_o0;
  wire  and2n_inst150_o0;
  wire  and2n_inst151_o0;
  wire  and2n_inst152_o0;
  wire  and2n_inst153_o0;
  wire  rr_func_cmpp_eq_inst15_0_stage_10_o0;
  wire  and2n_inst154_o0;
  wire  and2n_inst155_o0;
  wire  and2n_inst156_o0;
  wire  and2n_inst157_o0;
  wire  and2n_inst158_o0;
  wire  and2n_inst159_o0;
  wire  rr_func_cmpp_eq_inst16_stage_10_o0;
  wire  and2n_inst160_o0;
  wire  rr_func_cmpp_eq_inst16_stage_11_o0;
  wire  and2n_inst161_o0;
  wire  rr_func_cmpp_eq_inst16_stage_12_o0;
  wire  and2n_inst162_o0;
  wire  and2n_inst163_o0;
  wire  and2n_inst164_o0;
  wire  or3n_inst18_o0;
  wire  or3n_inst19_o0;
  wire  and2n_inst165_o0;
  wire  and2n_inst166_o0;
  wire  and2n_inst167_o0;
  wire  and2n_inst168_o0;
  wire  and2n_inst169_o0;
  wire  and2n_inst170_o0;
  wire  or2n_inst29_o0;
  wire  or3n_inst20_o0;
  wire  or2n_inst30_o0;
  wire  or2n_inst31_o0;
  wire  or3n_inst21_o0;
  wire  inverter1n_inst17_o0;
  wire  rr_func_cmpp_eq_inst17_stage_12_o0;
  wire  rr_func_cmpp_eq_inst17_0_stage_12_o0;
  wire [1 : 0] select_2_1_wn_inst9_o0;
  wire [1 : 0] select_2_1_wn_inst10_o0;
  wire  and2n_inst172_o0;
  wire [1 : 0] sext_inst74_o0;
  wire  or3n_inst22_o0;
  wire  or2n_inst34_o0;
  wire  and2n_inst174_o0;
  wire [1 : 0] rr_var_vactive_stage_13_o0;
  wire  and2n_inst171_o0;
  wire  inverter1n_inst18_o0;
  wire  or3n_inst23_o0;
  wire  or3n_inst24_o0;
  wire  or2n_inst35_o0;
  wire  and2n_inst173_o0;
  wire  inverter1n_inst19_o0;
  wire  and2n_inst175_o0;
  wire  and2n_inst176_o0;
  wire  and2n_inst177_o0;
  wire  and2n_inst178_o0;
  wire  and2n_inst179_o0;
  wire  and2n_inst180_o0;
  wire  and2n_inst181_o0;
  wire  and2n_inst182_o0;
  wire  and2n_inst183_o0;
  wire [31 : 0] rr_func_addw_inst8_stage_1_o0;
  wire  and2n_inst184_o0;
  wire  and2n_inst185_o0;
  wire  and2n_inst186_o0;
  wire  rr_func_cmpp_eq_inst18_stage_3_o0;
  wire  and2n_inst187_o0;
  wire  rr_func_cmpp_eq_inst18_stage_4_o0;
  wire  and2n_inst188_o0;
  wire  rr_func_cmpp_eq_inst18_stage_5_o0;
  wire  and2n_inst189_o0;
  wire  rr_func_cmpp_eq_inst18_stage_6_o0;
  wire  and2n_inst190_o0;
  wire  rr_func_cmpp_eq_inst18_stage_7_o0;
  wire  and2n_inst191_o0;
  wire  rr_func_cmpp_eq_inst18_stage_8_o0;
  wire  and2n_inst192_o0;
  wire  rr_func_cmpp_eq_inst18_stage_9_o0;
  wire  and2n_inst193_o0;
  wire  rr_func_cmpp_eq_inst18_stage_10_o0;
  wire  and2n_inst194_o0;
  wire  and2n_inst195_o0;
  wire  and2n_inst196_o0;
  wire  and2n_inst197_o0;
  wire  and2n_inst198_o0;
  wire  and2n_inst199_o0;
  wire  or3n_inst25_o0;
  wire  or2n_inst36_o0;
  wire  or3n_inst26_o0;
  wire  inverter1n_inst20_o0;
  wire [11 : 0] select_2_1_wn_inst11_o0;
  wire [11 : 0] select_2_1_wn_inst12_o0;
  wire  and2n_inst201_o0;
  wire [11 : 0] sext_inst75_o0;
  wire  and2n_inst203_o0;
  wire [11 : 0] rr_var_xa_stage_4_o0;
  wire  and2n_inst200_o0;
  wire  inverter1n_inst21_o0;
  wire  or3n_inst27_o0;
  wire  and2n_inst202_o0;
  wire  inverter1n_inst22_o0;
  wire  or3n_inst28_o0;
  wire  and2n_inst204_o0;
  wire  and2n_inst205_o0;
  wire  and2n_inst206_o0;
  wire  and2n_inst207_o0;
  wire  or2n_inst39_o0;
  wire  or3n_inst29_o0;
  wire  or3n_inst30_o0;
  wire  inverter1n_inst23_o0;
  wire [1 : 0] select_2_1_wn_inst13_o0;
  wire [1 : 0] select_2_1_wn_inst14_o0;
  wire  and2n_inst209_o0;
  wire  or2n_inst42_o0;
  wire  and2n_inst211_o0;
  wire  and2n_inst208_o0;
  wire  inverter1n_inst24_o0;
  wire  or3n_inst31_o0;
  wire  or2n_inst43_o0;
  wire  and2n_inst210_o0;
  wire  inverter1n_inst25_o0;
  wire  or3n_inst32_o0;
  wire  or2n_inst44_o0;
  wire  and2n_inst212_o0;
  wire  and2n_inst213_o0;
  wire  and2n_inst214_o0;
  wire  and2n_inst215_o0;
  wire  and2n_inst216_o0;
  wire  or2n_inst45_o0;
  wire  or3n_inst33_o0;
  wire  or2n_inst46_o0;
  wire  or3n_inst34_o0;
  wire  inverter1n_inst26_o0;
  wire [1 : 0] select_2_1_wn_inst15_o0;
  wire [1 : 0] select_2_1_wn_inst16_o0;
  wire  and2n_inst218_o0;
  wire  or3n_inst35_o0;
  wire  and2n_inst220_o0;
  wire  and2n_inst217_o0;
  wire  inverter1n_inst27_o0;
  wire  or3n_inst36_o0;
  wire  or2n_inst49_o0;
  wire  or2n_inst50_o0;
  wire  and2n_inst219_o0;
  wire  inverter1n_inst28_o0;
  wire  or3n_inst37_o0;
  wire  or2n_inst51_o0;
  wire  and2n_inst221_o0;
  wire  and2n_inst222_o0;
  wire  and2n_inst223_o0;
  wire  and2n_inst224_o0;
  wire  and2n_inst225_o0;
  wire  or2n_inst52_o0;
  wire  or3n_inst38_o0;
  wire  or2n_inst53_o0;
  wire  or3n_inst39_o0;
  wire  inverter1n_inst29_o0;
  wire [1 : 0] select_2_1_wn_inst17_o0;
  wire [1 : 0] select_2_1_wn_inst18_o0;
  wire  and2n_inst227_o0;
  wire  or3n_inst40_o0;
  wire  and2n_inst229_o0;
  wire  and2n_inst226_o0;
  wire  inverter1n_inst30_o0;
  wire  or3n_inst41_o0;
  wire  or2n_inst56_o0;
  wire  or2n_inst57_o0;
  wire  and2n_inst228_o0;
  wire  inverter1n_inst31_o0;
  wire  and2n_inst230_o0;
  wire  and2n_inst231_o0;
  wire  rr_func_cmpp_eq_inst22_stage_4_o0;
  wire  and2n_inst232_o0;
  wire  rr_func_cmpp_eq_inst22_stage_5_o0;
  wire  and2n_inst233_o0;
  wire  rr_func_cmpp_eq_inst22_stage_6_o0;
  wire  and2n_inst234_o0;
  wire  rr_func_cmpp_eq_inst22_stage_7_o0;
  wire  and2n_inst235_o0;
  wire  rr_func_cmpp_eq_inst22_stage_8_o0;
  wire  and2n_inst236_o0;
  wire  rr_func_cmpp_eq_inst22_stage_9_o0;
  wire  and2n_inst237_o0;
  wire  and2n_inst238_o0;
  wire  and2n_inst239_o0;
  wire  and2n_inst240_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_4_o0;
  wire  and2n_inst241_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_5_o0;
  wire  and2n_inst242_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_6_o0;
  wire  and2n_inst243_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_7_o0;
  wire  and2n_inst244_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_8_o0;
  wire  and2n_inst245_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_9_o0;
  wire  and2n_inst246_o0;
  wire  rr_func_cmpp_eq_inst22_0_stage_10_o0;
  wire  and2n_inst247_o0;
  wire  and2n_inst248_o0;
  wire  and2n_inst249_o0;
  wire  rr_func_cmpp_neq_inst0_stage_11_o0;
  wire  and2n_inst250_o0;
  wire  and2n_inst251_o0;
  wire  and2n_inst252_o0;
  wire  and2n_inst253_o0;
  wire  and2n_inst254_o0;
  wire  and2n_inst255_o0;
  wire  and2n_inst256_o0;
  wire [31 : 0] rr_func_addw_inst9_stage_5_o0;
  wire  and2n_inst257_o0;
  wire  and2n_inst258_o0;
  wire  and2n_inst259_o0;
  wire  rr_func_cmpp_eq_inst19_stage_7_o0;
  wire  and2n_inst260_o0;
  wire  rr_func_cmpp_eq_inst19_stage_8_o0;
  wire  and2n_inst261_o0;
  wire  rr_func_cmpp_eq_inst19_stage_9_o0;
  wire  and2n_inst262_o0;
  wire  rr_func_cmpp_eq_inst19_stage_10_o0;
  wire  and2n_inst263_o0;
  wire  rr_func_cmpp_eq_inst19_stage_11_o0;
  wire  and2n_inst264_o0;
  wire  and2n_inst265_o0;
  wire  or3n_inst42_o0;
  wire  or2n_inst58_o0;
  wire  and2n_inst266_o0;
  wire  and2n_inst267_o0;
  wire  and2n_inst268_o0;
  wire  and2n_inst269_o0;
  wire  and2n_inst270_o0;
  wire  or2n_inst59_o0;
  wire  or3n_inst43_o0;
  wire  or2n_inst60_o0;
  wire  or3n_inst44_o0;
  wire  inverter1n_inst32_o0;
  wire  rr_func_cmpp_eq_inst24_stage_10_o0;
  wire  rr_func_cmpp_eq_inst24_0_stage_10_o0;
  wire  rr_func_cmpp_eq_inst23_stage_10_o0;
  wire [1 : 0] select_2_1_wn_inst19_o0;
  wire [1 : 0] select_2_1_wn_inst20_o0;
  wire  and2n_inst272_o0;
  wire [1 : 0] sext_inst76_o0;
  wire  or3n_inst45_o0;
  wire  and2n_inst274_o0;
  wire [1 : 0] rr_var_cbarsactive_stage_11_o0;
  wire  and2n_inst271_o0;
  wire  inverter1n_inst33_o0;
  wire  or3n_inst46_o0;
  wire  or2n_inst63_o0;
  wire  or2n_inst64_o0;
  wire  and2n_inst273_o0;
  wire  inverter1n_inst34_o0;
  wire  and2n_inst275_o0;
  wire  and2n_inst276_o0;
  wire  or2n_inst65_o0;
  wire  or3n_inst47_o0;
  wire  inverter1n_inst35_o0;
  wire  rr_func_cmpp_eq_inst23_0_stage_10_o0;
  wire [1 : 0] select_2_1_wn_inst21_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst33_o0;
  wire  and2n_inst278_o0;
  wire  and2n_inst280_o0;
  wire [1 : 0] rr_var_castactive_stage_11_o0;
  wire  and2n_inst277_o0;
  wire  inverter1n_inst36_o0;
  wire  or2n_inst67_o0;
  wire  and3n_inst3_o0;
  wire  and2n_inst279_o0;
  wire  nor2n_inst2_o0;
  wire  nor2n_inst7_o0;
  wire  and2n_inst281_o0;
  wire  and2n_inst282_o0;
  wire  rr_func_cmpp_eq_inst23_stage_8_o0;
  wire  and2n_inst283_o0;
  wire  rr_func_cmpp_eq_inst23_stage_9_o0;
  wire  and2n_inst284_o0;
  wire  and2n_inst285_o0;
  wire  rr_func_cmpp_eq_inst23_stage_11_o0;
  wire  and2n_inst286_o0;
  wire  and2n_inst287_o0;
  wire  and2n_inst288_o0;
  wire  and2n_inst289_o0;
  wire  or3n_inst48_o0;
  wire  and2n_inst290_o0;
  wire  and2n_inst291_o0;
  wire  and2n_inst292_o0;
  wire  and2n_inst293_o0;
  wire  or2n_inst68_o0;
  wire  or3n_inst49_o0;
  wire  or3n_inst50_o0;
  wire  inverter1n_inst37_o0;
  wire  rr_func_cmpp_eq_inst20_0_stage_7_o0;
  wire  rr_func_cmpp_eq_inst21_stage_7_o0;
  wire  rr_func_cmpp_eq_inst21_0_stage_7_o0;
  wire [11 : 0] select_2_1_wn_inst22_o0;
  wire [11 : 0] select_2_1_wn_inst23_o0;
  wire  and2n_inst295_o0;
  wire  or2n_inst71_o0;
  wire  and2n_inst297_o0;
  wire  and2n_inst294_o0;
  wire  inverter1n_inst38_o0;
  wire  or3n_inst51_o0;
  wire  or2n_inst72_o0;
  wire  and2n_inst296_o0;
  wire  inverter1n_inst39_o0;
  wire  and2n_inst298_o0;
  wire [11 : 0] rr_var_ya_1_stage_9_o0;
  wire  and2n_inst299_o0;
  wire  and2n_inst300_o0;
  wire  and2n_inst301_o0;
  wire  and2n_inst302_o0;
  wire  and2n_inst303_o0;
  wire  and2n_inst304_o0;
  wire  and2n_inst305_o0;
  wire  and2n_inst306_o0;
  wire  and2n_inst307_o0;
  wire  and2n_inst308_o0;
  wire  and2n_inst309_o0;
  wire  and2n_inst310_o0;
  wire  rr_func_cmpp_neq_inst1_0_stage_11_o0;
  wire  and2n_inst311_o0;
  wire  and2n_inst312_o0;
  wire  and2n_inst313_o0;
  wire  and2n_inst314_o0;
  wire  and2n_inst315_o0;
  wire  and2n_inst316_o0;
  wire  and2n_inst317_o0;
  wire  rr_func_cmpp_eq_inst8_stage_12_o0;
  wire  and2n_inst318_o0;
  wire  and2n_inst319_o0;
  wire  and2n_inst320_o0;
  wire  and2n_inst321_o0;
  wire  and2n_inst322_o0;
  wire  and2n_inst323_o0;
  wire  and2n_inst324_o0;
  wire  and2n_inst325_o0;
  wire  and2n_inst326_o0;
  wire  and2n_inst327_o0;
  wire  and2n_inst328_o0;
  wire  and2n_inst329_o0;
  wire  and2n_inst330_o0;
  wire  and2n_inst331_o0;
  wire  and2n_inst332_o0;
  wire  and2n_inst333_o0;
  wire  and2n_inst334_o0;
  wire  and2n_inst335_o0;
  wire  and2n_inst336_o0;
  wire  rr_func_cmpp_eq_inst20_0_stage_3_o0;
  wire  and2n_inst337_o0;
  wire  rr_func_cmpp_eq_inst20_0_stage_4_o0;
  wire  and2n_inst338_o0;
  wire  rr_func_cmpp_eq_inst20_0_stage_5_o0;
  wire  and2n_inst339_o0;
  wire  and2n_inst340_o0;
  wire  and2n_inst341_o0;
  wire  and2n_inst342_o0;
  wire  and2n_inst343_o0;
  wire  and2n_inst344_o0;
  wire  and2n_inst345_o0;
  wire  and2n_inst346_o0;
  wire  and2n_inst347_o0;
  wire  and2n_inst348_o0;
  wire  and2n_inst349_o0;
  wire  and2n_inst350_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst24_o0;
  wire [1 : 0] sext_inst77_o0;
  wire [1 : 0] sext_inst78_o0;
  wire  or3n_inst53_o0;
  wire [1 : 0] sext_inst79_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst27_o0;
  wire [1 : 0] sext_inst80_o0;
  wire  nor2n_inst4_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst29_o0;
  wire [1 : 0] sext_inst81_o0;
  wire  or3n_inst56_o0;
  wire [1 : 0] sext_inst82_o0;
  wire [11 : 0] sext_inst83_o0;
  wire  inverter1n_inst40_o0;
  wire  or2n_inst80_o0;
  wire  or2n_inst81_o0;
  wire [11 : 0] sext_inst84_o0;
  wire  or2n_inst84_o0;
  wire [1 : 0] sext_inst85_o0;
  wire [1 : 0] sext_inst86_o0;
  wire  nor2n_inst6_o0;
  wire [1 : 0] sext_inst87_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst35_o0;
  wire [8 : 0] sext_inst88_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst37_o0;
  wire [8 : 0] sext_inst89_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst38_o0;
  wire [8 : 0] sext_inst90_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst39_o0;
  wire [8 : 0] sext_inst91_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst40_o0;
  wire [8 : 0] sext_inst92_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst42_o0;
  wire [8 : 0] sext_inst93_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst43_o0;
  wire [8 : 0] sext_inst94_o0;
  wire [8 : 0] datamerge_select_2_1_wn_inst44_o0;
  wire [8 : 0] sext_inst95_o0;
  wire [1 : 0] datamerge_select_2_1_wn_inst45_o0;
  wire  and2n_inst351_o0;
  wire  and2n_inst352_o0;
  wire  and2n_inst353_o0;
  wire  and2n_inst354_o0;
  wire  and2n_inst355_o0;
  wire  and2n_inst356_o0;
  wire  and2n_inst357_o0;
  wire  and2n_inst358_o0;
  wire  and2n_inst359_o0;
  wire  and2n_inst360_o0;
  wire  and2n_inst361_o0;
  wire  inverter1n_inst41_o0;
  wire  retimed_reg_o0;


  // Signal assignments

  assign err = 1'b0;
  assign sig_enable = enable;
  assign sig_start = start;
  assign sig_abort = abort;
  assign status = delayed_done_o0;
  assign sig_stallbar_in = stallbar_in;
  assign stallbar_out = inverter1n_inst42_o0;
  assign busy = or2n_inst2_o0;
  assign outstream_dvi_out_do_0 = outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_str_dataout;
  assign outstream_dvi_out_req_0 = outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_str_req;
  assign sig_outstream_dvi_out_ready_0 = outstream_dvi_out_ready_0;
  assign sig_lid_rawdatain_hsync_0_0 = lid_rawdatain_hsync_0_0;
  assign sig_lien_rawdatain_hsync_0_0 = lien_rawdatain_hsync_0_0;
  assign sig_lid_rawdatain_hblank_0_0 = lid_rawdatain_hblank_0_0;
  assign sig_lien_rawdatain_hblank_0_0 = lien_rawdatain_hblank_0_0;
  assign sig_lid_rawdatain_hbporch_0_0 = lid_rawdatain_hbporch_0_0;
  assign sig_lien_rawdatain_hbporch_0_0 = lien_rawdatain_hbporch_0_0;
  assign sig_lid_rawdatain_hactive_0_0 = lid_rawdatain_hactive_0_0;
  assign sig_lien_rawdatain_hactive_0_0 = lien_rawdatain_hactive_0_0;
  assign sig_lid_rawdatain_vsync_0_0 = lid_rawdatain_vsync_0_0;
  assign sig_lien_rawdatain_vsync_0_0 = lien_rawdatain_vsync_0_0;
  assign sig_lid_rawdatain_vblank_0_0 = lid_rawdatain_vblank_0_0;
  assign sig_lien_rawdatain_vblank_0_0 = lien_rawdatain_vblank_0_0;
  assign sig_lid_rawdatain_vbporch_0_0 = lid_rawdatain_vbporch_0_0;
  assign sig_lien_rawdatain_vbporch_0_0 = lien_rawdatain_vbporch_0_0;
  assign sig_lid_rawdatain_vactive_0_0 = lid_rawdatain_vactive_0_0;
  assign sig_lien_rawdatain_vactive_0_0 = lien_rawdatain_vactive_0_0;
  assign sig_lid_rawdatain_hfporch_0_0 = lid_rawdatain_hfporch_0_0;
  assign sig_lien_rawdatain_hfporch_0_0 = lien_rawdatain_hfporch_0_0;
  assign sig_lid_rawdatain_vfporch_0_0 = lid_rawdatain_vfporch_0_0;
  assign sig_lien_rawdatain_vfporch_0_0 = lien_rawdatain_vfporch_0_0;

  // Basic logic assignments


  // Component port and generic maps / Behavioural code.

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:117:28   Scheduled at time 8 (phase 0)
  mpylw_multi_stage_noreset #(.inwidth(0), .inwidth0(32), .inwidth1(2), .outwidth(32), .outlsb(0), .numstage(2))  mpylw_multi_stage_noreset_inst0(
                      .clk(clk),
                      .reset(reset),
                      .enable(and3n_inst0_o0),
                      .flush(1'b0),
                      .o0_enable(mpylw_multi_stage_noreset_inst0_o0_enable),
                      .pred(cmpp_eq_inst23_o1),
                      .i0(sr_var_vactive_1_o0[31 : 0]),
                      .i1(2'b11),
                      .o0(mpylw_multi_stage_noreset_inst0_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:139:3   Scheduled at time 13 (phase 0)
  test_pattern_generator_wide_ststream0_0_noreset #(.signwidth(6), .sdwidth(27), .strid(0), .dwidth0(8), .dwidth1(8), .dwidth2(8), .dwidth3(1), .dwidth4(1), .dwidth5(1))  outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0(
                      .clk(clk),
                      .reset(reset),
                      .enable(and3n_inst0_o0),
                      .flush(1'b0),
                      .str_ready(sig_outstream_dvi_out_ready_0),
                      .sign(outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_combine6_wn_inst0_o0[5 : 0]),
                      .str_req(outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_str_req),
                      .stallbar(outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_stallbar),
                      .pred(interconnect_select_1_1_wn_inst0_o0),
                      .str_dataout(outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_str_dataout[26 : 0]),
                      .datain0(datamerge_select_3_1_wn_inst10_o0[7 : 0]),
                      .datain1(datamerge_select_3_1_wn_inst11_o0[7 : 0]),
                      .datain2(datamerge_select_2_1_wn_inst41_o0[7 : 0]),
                      .datain3(rr_var_dvi_ds_s_hs_stage_12_o0),
                      .datain4(datamerge_select_3_1_wn_inst3_o0),
                      .datain5(datamerge_select_2_1_wn_inst45_o0[0]));

  brf #(.lcwidth(1))  brf_inst0(
                      .running(phasebus_0),
                      .enable(and3n_inst0_o0),
                      .p_enable(brf_inst0_p_enable),
                      .lc_enable(brf_inst0_lc_enable),
                      .op(1'b1),
                      .lc(sr_var_loopcounter_o0),
                      .p(brf_inst0_p),
                      .lc_out(brf_inst0_lc_out));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8   Scheduled at time 3 (phase 0)
  cmpp_eq_1 #(.width(12))  cmpp_eq_inst0(
                      .o0_enable(cmpp_eq_inst0_o0_enable),
                      .o1_enable(cmpp_eq_inst0_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_3_o0),
                      .i0(rr_var_x_stage_3_o0[11 : 0]),
                      .i1(sext_inst16_o0[11 : 0]),
                      .o0(cmpp_eq_inst0_o0),
                      .o1(cmpp_eq_inst0_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8   Scheduled at time 7 (phase 0)
  cmpp_eq_1 #(.width(12))  cmpp_eq_inst1(
                      .o0_enable(cmpp_eq_inst1_o0_enable),
                      .o1_enable(cmpp_eq_inst1_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_7_o0),
                      .i0(rr_var_y_stage_7_o0[11 : 0]),
                      .i1(sext_inst20_o0[11 : 0]),
                      .o0(cmpp_eq_inst1_o0),
                      .o1(cmpp_eq_inst1_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:107:7   Scheduled at time 4 (phase 0)   Speculated
  addw #(.width(12))  addw_inst0(
                      .o0_enable(addw_inst0_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_4_o0),
                      .i0(datamerge_select_2_1_wn_inst30_o0[11 : 0]),
                      .i1(sext_inst38_o0[11 : 0]),
                      .o0(addw_inst0_o0[11 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:145:6   Scheduled at time 7 (phase 0)   Speculated
  addw #(.width(12))  addw_inst1(
                      .o0_enable(addw_inst1_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_7_o0),
                      .i0(rr_var_y_stage_7_o0[11 : 0]),
                      .i1(sext_inst68_o0[11 : 0]),
                      .o0(addw_inst1_o0[11 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:146:8   Scheduled at time 8 (phase 0)   Speculated
  addw #(.width(12))  addw_inst2(
                      .o0_enable(addw_inst2_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_8_o0),
                      .i0(datamerge_select_2_1_wn_inst32_o0[11 : 0]),
                      .i1(sext_inst69_o0[11 : 0]),
                      .o0(addw_inst2_o0[11 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:150:5   Scheduled at time 3 (phase 0)   Speculated
  addw #(.width(12))  addw_inst3(
                      .o0_enable(addw_inst3_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_3_o0),
                      .i0(rr_var_x_stage_3_o0[11 : 0]),
                      .i1(sext_inst70_o0[11 : 0]),
                      .o0(addw_inst3_o0[11 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:73:24   Scheduled at time 7 (phase 0)
  cmpp_eq_1 #(.width(1))  cmpp_eq_inst2(
                      .o0_enable(cmpp_eq_inst2_o0_enable),
                      .o1_enable(cmpp_eq_inst2_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst0_stage_6_o0),
                      .i0(sr_var_hsync_o0),
                      .i1(1'b0),
                      .o0(cmpp_eq_inst2_o0),
                      .o1(cmpp_eq_inst2_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:75:24   Scheduled at time 7 (phase 0)
  cmpp_eq_1 #(.width(1))  cmpp_eq_inst3(
                      .o0_enable(cmpp_eq_inst3_o0_enable),
                      .o1_enable(cmpp_eq_inst3_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst12_stage_6_o0),
                      .i0(sr_var_hsync_o0),
                      .i1(1'b0),
                      .o0(cmpp_eq_inst3_o0),
                      .o1(cmpp_eq_inst3_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:83:24   Scheduled at time 13 (phase 0)
  cmpp_eq_1 #(.width(1))  cmpp_eq_inst4(
                      .o0_enable(cmpp_eq_inst4_o0_enable),
                      .o1_enable(cmpp_eq_inst4_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst1_stage_12_o0),
                      .i0(sr_var_vsync_o0),
                      .i1(1'b0),
                      .o0(cmpp_eq_inst4_o0),
                      .o1(cmpp_eq_inst4_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:85:24   Scheduled at time 13 (phase 0)
  cmpp_eq_1 #(.width(1))  cmpp_eq_inst5(
                      .o0_enable(cmpp_eq_inst5_o0_enable),
                      .o1_enable(cmpp_eq_inst5_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst15_stage_12_o0),
                      .i0(sr_var_vsync_o0),
                      .i1(1'b0),
                      .o0(cmpp_eq_inst5_o0),
                      .o1(cmpp_eq_inst5_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:8   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:104:15   Scheduled at time 11 (phase 0)   Speculated
  cmpr_neq #(.width(2))  cmpr_neq_inst0(
                      .o0_enable(cmpr_neq_inst0_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_11_o0),
                      .i0(interconnect_select_3_1_wn_inst0_o0[1 : 0]),
                      .i1(sext_inst35_o0[1 : 0]),
                      .o0(cmpr_neq_inst0_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:20   Scheduled at time 12 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst1(
                      .o0_enable(cmpr_neq_inst1_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_neq_inst0_0_stage_11_o0),
                      .i0(rr_var_ractive_stage_12_o0[1 : 0]),
                      .i1(sext_inst27_o0[1 : 0]),
                      .o0(cmpr_neq_inst1_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:99:16   Scheduled at time 12 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst2(
                      .o0_enable(cmpr_neq_inst2_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_12_o0),
                      .i0(rr_var_gactive_stage_12_o0[1 : 0]),
                      .i1(sext_inst30_o0[1 : 0]),
                      .o0(cmpr_neq_inst2_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:102:16   Scheduled at time 12 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst3(
                      .o0_enable(cmpr_neq_inst3_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_12_o0),
                      .i0(rr_var_ractive_stage_12_o0[1 : 0]),
                      .i1(sext_inst33_o0[1 : 0]),
                      .o0(cmpr_neq_inst3_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:19   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:125:19   Scheduled at time 13 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst4(
                      .o0_enable(cmpr_neq_inst4_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_neq_inst2_stage_12_o0),
                      .i0(rr_var_bactive_stage_12_o0[1 : 0]),
                      .i1(sext_inst43_o0[1 : 0]),
                      .o0(cmpr_neq_inst4_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:31   Scheduled at time 12 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst5(
                      .o0_enable(cmpr_neq_inst5_o0_enable),
                      .op(1'b0),
                      .pred(cmpp_eq_inst8_o1),
                      .i0(datamerge_select_3_1_wn_inst7_o0[1 : 0]),
                      .i1(sext_inst45_o0[1 : 0]),
                      .o0(cmpr_neq_inst5_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:125:31   Scheduled at time 12 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst6(
                      .o0_enable(cmpr_neq_inst6_o0_enable),
                      .op(1'b0),
                      .pred(cmpp_eq_inst8_o1),
                      .i0(datamerge_select_3_1_wn_inst6_o0[1 : 0]),
                      .i1(sext_inst49_o0[1 : 0]),
                      .o0(cmpr_neq_inst6_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:137:17   Scheduled at time 13 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst7(
                      .o0_enable(cmpr_neq_inst7_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_13_o0),
                      .i0(datamerge_select_3_1_wn_inst2_o0[1 : 0]),
                      .i1(sext_inst63_o0[1 : 0]),
                      .o0(cmpr_neq_inst7_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:137:28   Scheduled at time 13 (phase 0)
  cmpr_neq #(.width(2))  cmpr_neq_inst8(
                      .o0_enable(cmpr_neq_inst8_o0_enable),
                      .op(1'b0),
                      .pred(cmpp_eq_inst11_o1),
                      .i0(datamerge_select_3_1_wn_inst4_o0[1 : 0]),
                      .i1(sext_inst65_o0[1 : 0]),
                      .o0(cmpr_neq_inst8_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:7   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:104:14   Scheduled at time 11 (phase 0)   Speculated
  cmpr_eq #(.width(2))  cmpr_eq_inst0(
                      .o0_enable(cmpr_eq_inst0_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_11_o0),
                      .i0(cmpr_neq_inst0_o0[1 : 0]),
                      .i1(sext_inst36_o0[1 : 0]),
                      .o0(cmpr_eq_inst0_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:19   Scheduled at time 12 (phase 0)
  cmpr_eq #(.width(2))  cmpr_eq_inst1(
                      .o0_enable(cmpr_eq_inst1_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_neq_inst0_0_stage_11_o0),
                      .i0(cmpr_neq_inst1_o0[1 : 0]),
                      .i1(sext_inst28_o0[1 : 0]),
                      .o0(cmpr_eq_inst1_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:99:15   Scheduled at time 12 (phase 0)   Speculated
  cmpr_eq #(.width(2))  cmpr_eq_inst2(
                      .o0_enable(cmpr_eq_inst2_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_12_o0),
                      .i0(cmpr_neq_inst2_o0[1 : 0]),
                      .i1(sext_inst31_o0[1 : 0]),
                      .o0(cmpr_eq_inst2_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:102:15   Scheduled at time 12 (phase 0)   Speculated
  cmpr_eq #(.width(2))  cmpr_eq_inst3(
                      .o0_enable(cmpr_eq_inst3_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_brf_inst0_stage_12_o0),
                      .i0(cmpr_neq_inst3_o0[1 : 0]),
                      .i1(sext_inst34_o0[1 : 0]),
                      .o0(cmpr_eq_inst3_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:30   Scheduled at time 13 (phase 0)
  cmpr_eq #(.width(2))  cmpr_eq_inst4(
                      .o0_enable(cmpr_eq_inst4_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_eq_inst8_0_stage_12_o0),
                      .i0(rr_func_cmpr_neq_inst5_stage_12_o0[1 : 0]),
                      .i1(sext_inst46_o0[1 : 0]),
                      .o0(cmpr_eq_inst4_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:125:30   Scheduled at time 13 (phase 0)
  cmpr_eq #(.width(2))  cmpr_eq_inst5(
                      .o0_enable(cmpr_eq_inst5_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_eq_inst8_0_stage_12_o0),
                      .i0(rr_func_cmpr_neq_inst6_stage_12_o0[1 : 0]),
                      .i1(sext_inst50_o0[1 : 0]),
                      .o0(cmpr_eq_inst5_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:7   Scheduled at time 11 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst0(
                      .o0_enable(cmpp_neq_inst0_o0_enable),
                      .o1_enable(cmpp_neq_inst0_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst22_stage_10_o0),
                      .i0(cmpr_neq_inst0_o0[1 : 0]),
                      .i1(sext_inst37_o0[1 : 0]),
                      .o0(cmpp_neq_inst0_o0),
                      .o1(cmpp_neq_inst0_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:122:6   Scheduled at time 11 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst1(
                      .o0_enable(cmpp_neq_inst1_o0_enable),
                      .o1_enable(cmpp_neq_inst1_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_11_o0),
                      .i0(datamerge_select_3_1_wn_inst8_o0[1 : 0]),
                      .i1(sext_inst41_o0[1 : 0]),
                      .o0(cmpp_neq_inst1_o0),
                      .o1(cmpp_neq_inst1_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:123:7   Scheduled at time 12 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst2(
                      .o0_enable(cmpp_neq_inst2_o0_enable),
                      .o1_enable(cmpp_neq_inst2_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst1_stage_11_o0),
                      .i0(datamerge_select_3_1_wn_inst9_o0[1 : 0]),
                      .i1(sext_inst42_o0[1 : 0]),
                      .o0(cmpp_neq_inst2_o0),
                      .o1(cmpp_neq_inst2_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:127:18   Scheduled at time 13 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst3(
                      .o0_enable(cmpp_neq_inst3_o0_enable),
                      .o1_enable(cmpp_neq_inst3_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst2_0_stage_12_o0),
                      .i0(rr_var_ractive_stage_12_o0[1 : 0]),
                      .i1(sext_inst53_o0[1 : 0]),
                      .o0(cmpp_neq_inst3_o0),
                      .o1(cmpp_neq_inst3_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:128:18   Scheduled at time 13 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst4(
                      .o0_enable(cmpp_neq_inst4_o0_enable),
                      .o1_enable(cmpp_neq_inst4_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst2_0_stage_12_o0),
                      .i0(rr_var_gactive_stage_12_o0[1 : 0]),
                      .i1(sext_inst55_o0[1 : 0]),
                      .o0(cmpp_neq_inst4_o0),
                      .o1(cmpp_neq_inst4_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:130:17   Scheduled at time 13 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst5(
                      .o0_enable(cmpp_neq_inst5_o0_enable),
                      .o1_enable(cmpp_neq_inst5_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst1_stage_12_o0),
                      .i0(rr_var_bactive_stage_12_o0[1 : 0]),
                      .i1(sext_inst57_o0[1 : 0]),
                      .o0(cmpp_neq_inst5_o0),
                      .o1(cmpp_neq_inst5_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:132:17   Scheduled at time 13 (phase 0)
  cmpp_neq_1 #(.width(2))  cmpp_neq_inst6(
                      .o0_enable(cmpp_neq_inst6_o0_enable),
                      .o1_enable(cmpp_neq_inst6_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst1_0_stage_12_o0),
                      .i0(rr_var_gactive_stage_12_o0[1 : 0]),
                      .i1(sext_inst59_o0[1 : 0]),
                      .o0(cmpp_neq_inst6_o0),
                      .o1(cmpp_neq_inst6_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:16   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:19   Scheduled at time 12 (phase 0)
  cmpp_eq_1 #(.width(2))  cmpp_eq_inst6(
                      .o0_enable(cmpp_eq_inst6_o0_enable),
                      .o1_enable(cmpp_eq_inst6_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst22_stage_11_o0),
                      .i0(datamerge_select_2_1_wn_inst31_o0[1 : 0]),
                      .i1(sext_inst29_o0[1 : 0]),
                      .o0(cmpp_eq_inst6_o0),
                      .o1(cmpp_eq_inst6_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:101:7   Scheduled at time 12 (phase 0)
  cmpp_eq_1 #(.width(2))  cmpp_eq_inst7(
                      .o0_enable(cmpp_eq_inst7_o0_enable),
                      .o1_enable(cmpp_eq_inst7_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst22_stage_11_o0),
                      .i0(rr_var_bactive_stage_12_o0[1 : 0]),
                      .i1(sext_inst32_o0[1 : 0]),
                      .o0(cmpp_eq_inst7_o0),
                      .o1(cmpp_eq_inst7_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:19   Scheduled at time 12 (phase 0)
  cmpp_eq_1 #(.width(2))  cmpp_eq_inst8(
                      .o0_enable(cmpp_eq_inst8_o0_enable),
                      .o1_enable(cmpp_eq_inst8_o1_enable),
                      .op(3'b001),
                      .pred(cmpp_neq_inst2_o0),
                      .i0(datamerge_select_3_1_wn_inst5_o0[1 : 0]),
                      .i1(sext_inst44_o0[1 : 0]),
                      .o0(cmpp_eq_inst8_o0),
                      .o1(cmpp_eq_inst8_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:27   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:30   Scheduled at time 13 (phase 0)
  cmpp_eq_1 #(.width(2))  cmpp_eq_inst9(
                      .o0_enable(cmpp_eq_inst9_o0_enable),
                      .o1_enable(cmpp_eq_inst9_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst2_stage_12_o0),
                      .i0(datamerge_select_2_1_wn_inst34_o0[1 : 0]),
                      .i1(sext_inst47_o0[1 : 0]),
                      .o0(cmpp_eq_inst9_o0),
                      .o1(cmpp_eq_inst9_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:125:27   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:125:30   Scheduled at time 13 (phase 0)
  cmpp_eq_1 #(.width(2))  cmpp_eq_inst10(
                      .o0_enable(cmpp_eq_inst10_o0_enable),
                      .o1_enable(cmpp_eq_inst10_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_neq_inst2_stage_12_o0),
                      .i0(datamerge_select_2_1_wn_inst36_o0[1 : 0]),
                      .i1(sext_inst51_o0[1 : 0]),
                      .o0(cmpp_eq_inst10_o0),
                      .o1(cmpp_eq_inst10_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:137:17   Scheduled at time 13 (phase 0)
  cmpp_eq_1 #(.width(2))  cmpp_eq_inst11(
                      .o0_enable(cmpp_eq_inst11_o0_enable),
                      .o1_enable(cmpp_eq_inst11_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_13_o0),
                      .i0(datamerge_select_3_1_wn_inst2_o0[1 : 0]),
                      .i1(sext_inst64_o0[1 : 0]),
                      .o0(cmpp_eq_inst11_o0),
                      .o1(cmpp_eq_inst11_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15   Scheduled at time 4 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst12(
                      .o0_enable(cmpp_eq_inst12_o0_enable),
                      .o1_enable(cmpp_eq_inst12_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst0_0_stage_3_o0),
                      .i0(sext_inst4_o0[31 : 0]),
                      .i1(sr_var_hblank_o0[31 : 0]),
                      .o0(cmpp_eq_inst12_o0),
                      .o1(cmpp_eq_inst12_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15   Scheduled at time 6 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst13(
                      .o0_enable(cmpp_eq_inst13_o0_enable),
                      .o1_enable(cmpp_eq_inst13_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst12_0_stage_5_o0),
                      .i0(sext_inst3_o0[31 : 0]),
                      .i1(rr_func_addw_inst4_stage_5_o0[31 : 0]),
                      .o0(cmpp_eq_inst13_o0),
                      .o1(cmpp_eq_inst13_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15   Scheduled at time 8 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst14(
                      .o0_enable(cmpp_eq_inst14_o0_enable),
                      .o1_enable(cmpp_eq_inst14_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst13_0_stage_7_o0),
                      .i0(sext_inst2_o0[31 : 0]),
                      .i1(rr_func_addw_inst5_stage_7_o0[31 : 0]),
                      .o0(cmpp_eq_inst14_o0),
                      .o1(cmpp_eq_inst14_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15   Scheduled at time 8 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst15(
                      .o0_enable(cmpp_eq_inst15_o0_enable),
                      .o1_enable(cmpp_eq_inst15_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst1_0_stage_7_o0),
                      .i0(sext_inst9_o0[31 : 0]),
                      .i1(sr_var_vblank_o0[31 : 0]),
                      .o0(cmpp_eq_inst15_o0),
                      .o1(cmpp_eq_inst15_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:15   Scheduled at time 10 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst16(
                      .o0_enable(cmpp_eq_inst16_o0_enable),
                      .o1_enable(cmpp_eq_inst16_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst15_0_stage_9_o0),
                      .i0(sext_inst8_o0[31 : 0]),
                      .i1(rr_func_addw_inst6_stage_9_o0[31 : 0]),
                      .o0(cmpp_eq_inst16_o0),
                      .o1(cmpp_eq_inst16_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:15   Scheduled at time 12 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst17(
                      .o0_enable(cmpp_eq_inst17_o0_enable),
                      .o1_enable(cmpp_eq_inst17_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst16_0_stage_11_o0),
                      .i0(sext_inst7_o0[31 : 0]),
                      .i1(rr_func_addw_inst7_stage_11_o0[31 : 0]),
                      .o0(cmpp_eq_inst17_o0),
                      .o1(cmpp_eq_inst17_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8   Scheduled at time 3 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst18(
                      .o0_enable(cmpp_eq_inst18_o0_enable),
                      .o1_enable(cmpp_eq_inst18_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_3_o0),
                      .i0(sext_inst1_o0[31 : 0]),
                      .i1(rr_func_addw_inst8_stage_2_o0[31 : 0]),
                      .o0(cmpp_eq_inst18_o0),
                      .o1(cmpp_eq_inst18_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8   Scheduled at time 7 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst19(
                      .o0_enable(cmpp_eq_inst19_o0_enable),
                      .o1_enable(cmpp_eq_inst19_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_7_o0),
                      .i0(sext_inst6_o0[31 : 0]),
                      .i1(rr_func_addw_inst9_stage_6_o0[31 : 0]),
                      .o0(cmpp_eq_inst19_o0),
                      .o1(cmpp_eq_inst19_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8   Scheduled at time 3 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst20(
                      .o0_enable(cmpp_eq_inst20_o0_enable),
                      .o1_enable(cmpp_eq_inst20_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_brf_inst0_stage_3_o0),
                      .i0(sext_inst0_o0[31 : 0]),
                      .i1(rr_func_addsubw_inst0_stage_2_o0[31 : 0]),
                      .o0(cmpp_eq_inst20_o0),
                      .o1(cmpp_eq_inst20_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:9   Scheduled at time 7 (phase 0)
  cmpp_eq_1 #(.width(32))  cmpp_eq_inst21(
                      .o0_enable(cmpp_eq_inst21_o0_enable),
                      .o1_enable(cmpp_eq_inst21_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst20_stage_6_o0),
                      .i0(sext_inst5_o0[31 : 0]),
                      .i1(rr_func_addsubw_inst1_stage_6_o0[31 : 0]),
                      .o0(cmpp_eq_inst21_o0),
                      .o1(cmpp_eq_inst21_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:25   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:25   Scheduled at time 5 (phase 0)
  addw #(.width(32))  addw_inst4(
                      .o0_enable(addw_inst4_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_cmpp_eq_inst12_0_stage_4_o0),
                      .i0(sr_var_hblank_o0[31 : 0]),
                      .i1(sr_var_hbporch_o0[31 : 0]),
                      .o0(addw_inst4_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:35   Scheduled at time 7 (phase 0)
  addw #(.width(32))  addw_inst5(
                      .o0_enable(addw_inst5_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_cmpp_eq_inst13_0_stage_6_o0),
                      .i0(rr_func_addw_inst4_stage_6_o0[31 : 0]),
                      .i1(sr_var_hactive_1_o0[31 : 0]),
                      .o0(addw_inst5_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:25   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:25   Scheduled at time 9 (phase 0)
  addw #(.width(32))  addw_inst6(
                      .o0_enable(addw_inst6_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_cmpp_eq_inst15_0_stage_8_o0),
                      .i0(sr_var_vblank_o0[31 : 0]),
                      .i1(sr_var_vbporch_o0[31 : 0]),
                      .o0(addw_inst6_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:35   Scheduled at time 11 (phase 0)
  addw #(.width(32))  addw_inst7(
                      .o0_enable(addw_inst7_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_cmpp_eq_inst16_0_stage_10_o0),
                      .i0(rr_func_addw_inst6_stage_10_o0[31 : 0]),
                      .i1(sr_var_vactive_1_o0[31 : 0]),
                      .o0(addw_inst7_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:18   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:28   Scheduled at time 0 (phase 0)
  addw #(.width(32))  addw_inst8(
                      .o0_enable(addw_inst8_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_0_o0),
                      .i0(sr_var_hblank_o0[31 : 0]),
                      .i1(sr_var_hbporch_o0[31 : 0]),
                      .o0(addw_inst8_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:18   dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:29   Scheduled at time 4 (phase 0)
  addw #(.width(32))  addw_inst9(
                      .o0_enable(addw_inst9_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_4_o0),
                      .i0(sr_var_vblank_o0[31 : 0]),
                      .i1(sr_var_vbporch_o0[31 : 0]),
                      .o0(addw_inst9_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:18   Scheduled at time 0 (phase 0)
  addw #(.width(32))  addw_inst10(
                      .o0_enable(addw_inst10_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_0_o0),
                      .i0(sr_var_hactive_1_o0[31 : 0]),
                      .i1(sr_var_hfporch_o0[31 : 0]),
                      .o0(addw_inst10_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:38   Scheduled at time 1 (phase 0)
  addw #(.width(32))  addw_inst11(
                      .o0_enable(addw_inst11_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_brf_inst0_stage_1_o0),
                      .i0(rr_func_addw_inst8_stage_0_o0[31 : 0]),
                      .i1(rr_func_addw_inst10_stage_0_o0[31 : 0]),
                      .o0(addw_inst11_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:19   Scheduled at time 4 (phase 0)
  addw #(.width(32))  addw_inst12(
                      .o0_enable(addw_inst12_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_cmpp_eq_inst20_stage_3_o0),
                      .i0(sr_var_vactive_1_o0[31 : 0]),
                      .i1(sr_var_vfporch_o0[31 : 0]),
                      .o0(addw_inst12_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:39   Scheduled at time 5 (phase 0)
  addw #(.width(32))  addw_inst13(
                      .o0_enable(addw_inst13_o0_enable),
                      .op(1'b1),
                      .pred(rr_func_cmpp_eq_inst20_stage_4_o0),
                      .i0(rr_func_addw_inst9_stage_4_o0[31 : 0]),
                      .i1(rr_func_addw_inst12_stage_4_o0[31 : 0]),
                      .o0(addw_inst13_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:48   Scheduled at time 2 (phase 0)
  addsubw #(.width(32))  addsubw_inst0(
                      .o0_enable(addsubw_inst0_o0_enable),
                      .op(2'b01),
                      .pred(rr_func_brf_inst0_stage_2_o0),
                      .i0(rr_func_addw_inst11_stage_1_o0[31 : 0]),
                      .i1(sext_inst66_o0[31 : 0]),
                      .o0(addsubw_inst0_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:49   Scheduled at time 6 (phase 0)
  addsubw #(.width(32))  addsubw_inst1(
                      .o0_enable(addsubw_inst1_o0_enable),
                      .op(2'b01),
                      .pred(rr_func_cmpp_eq_inst20_stage_5_o0),
                      .i0(rr_func_addw_inst13_stage_5_o0[31 : 0]),
                      .i1(sext_inst67_o0[31 : 0]),
                      .o0(addsubw_inst1_o0[31 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:26   Scheduled at time 4 (phase 0)
  shrkw #(.width(33), .shiftbits(3))  shrkw_inst0(
                      .o0_enable(shrkw_inst0_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_eq_inst18_0_stage_3_o0),
                      .i0(sext_inst14_o0[32 : 0]),
                      .o0(shrkw_inst0_o0[32 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:20   Scheduled at time 8 (phase 0)
  shrkw #(.width(33), .shiftbits(1))  shrkw_inst1(
                      .o0_enable(shrkw_inst1_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_eq_inst19_0_stage_7_o0),
                      .i0(sext_inst15_o0[32 : 0]),
                      .o0(shrkw_inst1_o0[32 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:117:31   Scheduled at time 9 (phase 0)
  shrkw #(.width(33), .shiftbits(2))  shrkw_inst2(
                      .o0_enable(shrkw_inst2_o0_enable),
                      .op(1'b0),
                      .pred(rr_func_cmpp_eq_inst23_0_stage_8_o0),
                      .i0(sext_inst13_o0[32 : 0]),
                      .o0(shrkw_inst2_o0[32 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16   Scheduled at time 4 (phase 0)
  cmpp_eq_1 #(.width(29))  cmpp_eq_inst22(
                      .o0_enable(cmpp_eq_inst22_o0_enable),
                      .o1_enable(cmpp_eq_inst22_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst18_0_stage_3_o0),
                      .i0(sext_inst10_o0[28 : 0]),
                      .i1(shrkw_inst0_o0[28 : 0]),
                      .o0(cmpp_eq_inst22_o0),
                      .o1(cmpp_eq_inst22_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10   Scheduled at time 8 (phase 0)
  cmpp_eq_1 #(.width(31))  cmpp_eq_inst23(
                      .o0_enable(cmpp_eq_inst23_o0_enable),
                      .o1_enable(cmpp_eq_inst23_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst19_0_stage_7_o0),
                      .i0(sext_inst12_o0[30 : 0]),
                      .i1(shrkw_inst1_o0[30 : 0]),
                      .o0(cmpp_eq_inst23_o0),
                      .o1(cmpp_eq_inst23_o1));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:117:17   Scheduled at time 10 (phase 0)
  cmpp_eq_1 #(.width(30))  cmpp_eq_inst24(
                      .o0_enable(cmpp_eq_inst24_o0_enable),
                      .o1_enable(cmpp_eq_inst24_o1_enable),
                      .op(3'b001),
                      .pred(rr_func_cmpp_eq_inst23_0_stage_9_o0),
                      .i0(sext_inst11_o0[29 : 0]),
                      .i1(rr_func_shrkw_inst2_stage_9_o0[29 : 0]),
                      .o0(cmpp_eq_inst24_o0),
                      .o1(cmpp_eq_inst24_o1));

  assign and3n_inst0_o0 = sig_enable & sig_stallbar_in & inverter1n_inst42_o0;

  sregn_noinit #(.width(1))  delayed_start(
                      .clk(clk),
                      .reset(reset),
                      .enable(and3n_inst0_o0),
                      .i0(sig_start),
                      .o0(startbus));

  rsflipflop_noinit  controller_rsflipflop_noinit_inst0(
                      .clk(clk),
                      .reset(reset),
                      .r(and2n_inst0_o0),
                      .s(and2n_inst2_o0),
                      .q(controller_rsflipflop_noinit_inst0_q));

  assign and2n_inst0_o0 = stagereg13_o0 & and3n_inst0_o0;
  assign inverter1n_inst0_o0 = ~and2n_inst0_o0;
  assign and2n_inst1_o0 = startbus & inverter1n_inst0_o0;
  assign and2n_inst2_o0 = and2n_inst1_o0 & and3n_inst0_o0;
  assign phasebus_0 = startbus | controller_rsflipflop_noinit_inst0_q;
  assign or2n_inst1_o0 = startbus | controller_rsflipflop_noinit_inst1_q;
  assign and2n_inst3_o0 = and2n_inst8_o0 & or2n_inst1_o0;

  rsflipflop_noinit  controller_rsflipflop_noinit_inst1(
                      .clk(clk),
                      .reset(reset),
                      .r(and2n_inst4_o0),
                      .s(and2n_inst6_o0),
                      .q(controller_rsflipflop_noinit_inst1_q));

  assign and2n_inst4_o0 = and2n_inst3_o0 & and3n_inst0_o0;
  assign and2n_inst5_o0 = startbus & and3n_inst0_o0;
  assign inverter1n_inst1_o0 = ~and2n_inst4_o0;
  assign and2n_inst6_o0 = inverter1n_inst1_o0 & and2n_inst5_o0;
  assign and2n_inst7_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  stagereg1(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(and2n_inst3_o0),
                      .o0(stagereg1_o0));

  sregn_noinit #(.width(1))  stagereg2(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg1_o0),
                      .o0(stagereg2_o0));

  sregn_noinit #(.width(1))  stagereg3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg2_o0),
                      .o0(stagereg3_o0));

  sregn_noinit #(.width(1))  stagereg4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg3_o0),
                      .o0(stagereg4_o0));

  sregn_noinit #(.width(1))  stagereg5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg4_o0),
                      .o0(stagereg5_o0));

  sregn_noinit #(.width(1))  stagereg6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg5_o0),
                      .o0(stagereg6_o0));

  sregn_noinit #(.width(1))  stagereg7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg6_o0),
                      .o0(stagereg7_o0));

  sregn_noinit #(.width(1))  stagereg8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg7_o0),
                      .o0(stagereg8_o0));

  sregn_noinit #(.width(1))  stagereg9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg8_o0),
                      .o0(stagereg9_o0));

  sregn_noinit #(.width(1))  stagereg10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg9_o0),
                      .o0(stagereg10_o0));

  sregn_noinit #(.width(1))  stagereg11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg10_o0),
                      .o0(stagereg11_o0));

  sregn_noinit #(.width(1))  stagereg12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg11_o0),
                      .o0(stagereg12_o0));

  sregn_noinit #(.width(1))  stagereg13(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst7_o0),
                      .i0(stagereg12_o0),
                      .o0(stagereg13_o0));

  sregn_noinit #(.width(1))  delayed_done(
                      .clk(clk),
                      .reset(reset),
                      .enable(and3n_inst0_o0),
                      .i0(stagereg13_o0),
                      .o0(delayed_done_o0));

  assign or2n_inst2_o0 = phasebus_0 | delayed_done_o0;

  combine6_wn #(.inwidth(1))  outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_combine6_wn_inst0(
                      .i0(1'b0),
                      .i1(1'b0),
                      .i2(1'b0),
                      .i3(1'b0),
                      .i4(1'b0),
                      .i5(1'b0),
                      .o0(outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_combine6_wn_inst0_o0[5 : 0]));

  assign and2n_inst8_o0 = phasebus_0 & equal_inst0_o0;

  equal #(.width(1))  equal_inst0(
                      .i0(sr_var_loopcounter_o0),
                      .i1(1'b0),
                      .o0(equal_inst0_o0));

  select_1_1_wn #(.dwidth(1))  interconnect_select_1_1_wn_inst0(
                      .enable0(phasebus_0),
                      .i0(rr_func_brf_inst0_stage_13_o0),
                      .o0(interconnect_select_1_1_wn_inst0_o0));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst0(
                      .i0(rr_var_x_stage_3_o0[11 : 0]),
                      .o0(sext_inst0_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst1(
                      .i0(rr_var_x_stage_3_o0[11 : 0]),
                      .o0(sext_inst1_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst2(
                      .i0(rr_var_x_stage_8_o0[11 : 0]),
                      .o0(sext_inst2_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst3(
                      .i0(rr_var_x_stage_6_o0[11 : 0]),
                      .o0(sext_inst3_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst4(
                      .i0(rr_var_x_stage_4_o0[11 : 0]),
                      .o0(sext_inst4_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst5(
                      .i0(rr_var_y_stage_7_o0[11 : 0]),
                      .o0(sext_inst5_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst6(
                      .i0(rr_var_y_stage_7_o0[11 : 0]),
                      .o0(sext_inst6_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst7(
                      .i0(rr_var_y_stage_12_o0[11 : 0]),
                      .o0(sext_inst7_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst8(
                      .i0(rr_var_y_stage_10_o0[11 : 0]),
                      .o0(sext_inst8_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(32), .signedflag(0))  sext_inst9(
                      .i0(rr_var_y_stage_8_o0[11 : 0]),
                      .o0(sext_inst9_o0[31 : 0]));

  sext #(.inwidth(12), .outwidth(29), .signedflag(0))  sext_inst10(
                      .i0(datamerge_select_2_1_wn_inst30_o0[11 : 0]),
                      .o0(sext_inst10_o0[28 : 0]));

  select_3_1_wn #(.dwidth(2))  interconnect_select_3_1_wn_inst0(
                      .enable0(rr_func_cmpp_eq_inst18_stage_11_o0),
                      .enable1(or2n_inst3_o0),
                      .enable2(rr_func_cmpp_eq_inst22_stage_11_o0),
                      .i0(sext_inst24_o0[1 : 0]),
                      .i1(rr_var_bactive_stage_12_o0[1 : 0]),
                      .i2(rr_func_moveii_inst40_stage_11_o0[1 : 0]),
                      .o0(interconnect_select_3_1_wn_inst0_o0[1 : 0]));

  assign or2n_inst3_o0 = rr_func_cmpp_eq_inst22_0_stage_11_o0 | nor3n_inst0_o0;

  sext #(.inwidth(12), .outwidth(30), .signedflag(0))  sext_inst11(
                      .i0(rr_var_ya_1_stage_10_o0[11 : 0]),
                      .o0(sext_inst11_o0[29 : 0]));

  sext #(.inwidth(12), .outwidth(31), .signedflag(0))  sext_inst12(
                      .i0(rr_var_ya_1_stage_8_o0[11 : 0]),
                      .o0(sext_inst12_o0[30 : 0]));

  sext #(.inwidth(32), .outwidth(33), .signedflag(0))  sext_inst13(
                      .i0(mpylw_multi_stage_noreset_inst0_o0[31 : 0]),
                      .o0(sext_inst13_o0[32 : 0]));

  sext #(.inwidth(32), .outwidth(33), .signedflag(0))  sext_inst14(
                      .i0(sr_var_hactive_1_o0[31 : 0]),
                      .o0(sext_inst14_o0[32 : 0]));

  sext #(.inwidth(32), .outwidth(33), .signedflag(0))  sext_inst15(
                      .i0(sr_var_vactive_1_o0[31 : 0]),
                      .o0(sext_inst15_o0[32 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst16(
                      .i0(1'b0),
                      .o0(sext_inst16_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst17(
                      .i0(1'b1),
                      .o0(sext_inst17_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst18(
                      .i0(1'b1),
                      .o0(sext_inst18_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst19(
                      .i0(1'b1),
                      .o0(sext_inst19_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst20(
                      .i0(1'b0),
                      .o0(sext_inst20_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst21(
                      .i0(1'b1),
                      .o0(sext_inst21_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst22(
                      .i0(1'b1),
                      .o0(sext_inst22_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst23(
                      .i0(1'b1),
                      .o0(sext_inst23_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst24(
                      .i0(1'b1),
                      .o0(sext_inst24_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst25(
                      .i0(1'b1),
                      .o0(sext_inst25_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst26(
                      .i0(1'b1),
                      .o0(sext_inst26_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst27(
                      .i0(1'b0),
                      .o0(sext_inst27_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst28(
                      .i0(1'b0),
                      .o0(sext_inst28_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst29(
                      .i0(1'b1),
                      .o0(sext_inst29_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst30(
                      .i0(1'b0),
                      .o0(sext_inst30_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst31(
                      .i0(1'b0),
                      .o0(sext_inst31_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst32(
                      .i0(1'b0),
                      .o0(sext_inst32_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst33(
                      .i0(1'b0),
                      .o0(sext_inst33_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst34(
                      .i0(1'b0),
                      .o0(sext_inst34_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst35(
                      .i0(1'b0),
                      .o0(sext_inst35_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst36(
                      .i0(1'b0),
                      .o0(sext_inst36_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst37(
                      .i0(1'b0),
                      .o0(sext_inst37_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst38(
                      .i0(1'b1),
                      .o0(sext_inst38_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst39(
                      .i0(1'b1),
                      .o0(sext_inst39_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst40(
                      .i0(1'b1),
                      .o0(sext_inst40_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst41(
                      .i0(1'b0),
                      .o0(sext_inst41_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst42(
                      .i0(1'b0),
                      .o0(sext_inst42_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst43(
                      .i0(1'b0),
                      .o0(sext_inst43_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst44(
                      .i0(1'b0),
                      .o0(sext_inst44_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst45(
                      .i0(1'b0),
                      .o0(sext_inst45_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst46(
                      .i0(1'b0),
                      .o0(sext_inst46_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst47(
                      .i0(1'b1),
                      .o0(sext_inst47_o0[1 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst48(
                      .i0(8'b11000000),
                      .o0(sext_inst48_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst49(
                      .i0(1'b0),
                      .o0(sext_inst49_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst50(
                      .i0(1'b0),
                      .o0(sext_inst50_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst51(
                      .i0(1'b1),
                      .o0(sext_inst51_o0[1 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst52(
                      .i0(8'b11000000),
                      .o0(sext_inst52_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst53(
                      .i0(1'b0),
                      .o0(sext_inst53_o0[1 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst54(
                      .i0(8'b11000000),
                      .o0(sext_inst54_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst55(
                      .i0(1'b0),
                      .o0(sext_inst55_o0[1 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst56(
                      .i0(8'b11000000),
                      .o0(sext_inst56_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst57(
                      .i0(1'b0),
                      .o0(sext_inst57_o0[1 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst58(
                      .i0(8'b11000000),
                      .o0(sext_inst58_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst59(
                      .i0(1'b0),
                      .o0(sext_inst59_o0[1 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst60(
                      .i0(8'b11111111),
                      .o0(sext_inst60_o0[8 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst61(
                      .i0(8'b11111111),
                      .o0(sext_inst61_o0[8 : 0]));

  sext #(.inwidth(8), .outwidth(9), .signedflag(0))  sext_inst62(
                      .i0(8'b11111111),
                      .o0(sext_inst62_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst63(
                      .i0(1'b0),
                      .o0(sext_inst63_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst64(
                      .i0(1'b0),
                      .o0(sext_inst64_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(0))  sext_inst65(
                      .i0(1'b0),
                      .o0(sext_inst65_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(32), .signedflag(0))  sext_inst66(
                      .i0(1'b1),
                      .o0(sext_inst66_o0[31 : 0]));

  sext #(.inwidth(1), .outwidth(32), .signedflag(0))  sext_inst67(
                      .i0(1'b1),
                      .o0(sext_inst67_o0[31 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst68(
                      .i0(1'b1),
                      .o0(sext_inst68_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst69(
                      .i0(1'b1),
                      .o0(sext_inst69_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst70(
                      .i0(1'b1),
                      .o0(sext_inst70_o0[11 : 0]));

  assign or2n_inst4_o0 = and2n_inst9_o0 | sig_start;
  assign and2n_inst9_o0 = brf_inst0_p_enable & phasebus_0;

  select_2_1_wn #(.dwidth(1))  select_2_1_wn_inst0(
                      .enable0(and2n_inst9_o0),
                      .enable1(and2n_inst11_o0),
                      .i0(brf_inst0_p),
                      .i1(1'b1),
                      .o0(select_2_1_wn_inst0_o0));

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_0(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst10_o0),
                      .i0(select_2_1_wn_inst0_o0),
                      .o0(rr_func_brf_inst0_stage_0_o0));

  assign and2n_inst10_o0 = or2n_inst4_o0 & and3n_inst0_o0;
  assign inverter1n_inst2_o0 = ~and2n_inst9_o0;
  assign and2n_inst11_o0 = sig_start & inverter1n_inst2_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_1(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst12_o0),
                      .i0(rr_func_brf_inst0_stage_0_o0),
                      .o0(rr_func_brf_inst0_stage_1_o0));

  assign and2n_inst12_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_2(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst13_o0),
                      .i0(rr_func_brf_inst0_stage_1_o0),
                      .o0(rr_func_brf_inst0_stage_2_o0));

  assign and2n_inst13_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst14_o0),
                      .i0(rr_func_brf_inst0_stage_2_o0),
                      .o0(rr_func_brf_inst0_stage_3_o0));

  assign and2n_inst14_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst15_o0),
                      .i0(rr_func_brf_inst0_stage_3_o0),
                      .o0(rr_func_brf_inst0_stage_4_o0));

  assign and2n_inst15_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst16_o0),
                      .i0(rr_func_brf_inst0_stage_4_o0),
                      .o0(rr_func_brf_inst0_stage_5_o0));

  assign and2n_inst16_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst17_o0),
                      .i0(rr_func_brf_inst0_stage_5_o0),
                      .o0(rr_func_brf_inst0_stage_6_o0));

  assign and2n_inst17_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst18_o0),
                      .i0(rr_func_brf_inst0_stage_6_o0),
                      .o0(rr_func_brf_inst0_stage_7_o0));

  assign and2n_inst18_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst19_o0),
                      .i0(rr_func_brf_inst0_stage_7_o0),
                      .o0(rr_func_brf_inst0_stage_8_o0));

  assign and2n_inst19_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst20_o0),
                      .i0(rr_func_brf_inst0_stage_8_o0),
                      .o0(rr_func_brf_inst0_stage_9_o0));

  assign and2n_inst20_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst21_o0),
                      .i0(rr_func_brf_inst0_stage_9_o0),
                      .o0(rr_func_brf_inst0_stage_10_o0));

  assign and2n_inst21_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst22_o0),
                      .i0(rr_func_brf_inst0_stage_10_o0),
                      .o0(rr_func_brf_inst0_stage_11_o0));

  assign and2n_inst22_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst23_o0),
                      .i0(rr_func_brf_inst0_stage_11_o0),
                      .o0(rr_func_brf_inst0_stage_12_o0));

  assign and2n_inst23_o0 = phasebus_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  rr_func_brf_inst0_stage_13(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst24_o0),
                      .i0(rr_func_brf_inst0_stage_12_o0),
                      .o0(rr_func_brf_inst0_stage_13_o0));

  assign and2n_inst24_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst25_o0 = cmpp_eq_inst0_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst26_o0),
                      .i0(cmpp_eq_inst0_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_3_o0));

  assign and2n_inst26_o0 = and2n_inst25_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst27_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_3_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_4_o0));

  assign and2n_inst27_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst28_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_5_o0));

  assign and2n_inst28_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst29_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_6_o0));

  assign and2n_inst29_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst30_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_7_o0));

  assign and2n_inst30_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst31_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_8_o0));

  assign and2n_inst31_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst32_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_9_o0));

  assign and2n_inst32_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst33_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_10_o0));

  assign and2n_inst33_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst34_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_11_o0));

  assign and2n_inst34_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst35_o0),
                      .i0(rr_func_cmpp_eq_inst0_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst0_stage_12_o0));

  assign and2n_inst35_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst36_o0 = cmpp_eq_inst0_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:72:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst0_0_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst37_o0),
                      .i0(cmpp_eq_inst0_o1),
                      .o0(rr_func_cmpp_eq_inst0_0_stage_3_o0));

  assign and2n_inst37_o0 = and2n_inst36_o0 & and3n_inst0_o0;
  assign or3n_inst1_o0 = and2n_inst38_o0 | and2n_inst39_o0 | and2n_inst40_o0;
  assign or2n_inst6_o0 = and2n_inst40_o0 | and2n_inst39_o0;
  assign or3n_inst2_o0 = or2n_inst6_o0 | sig_start | phasebus_0;
  assign inverter1n_inst3_o0 = ~or2n_inst6_o0;
  assign and2n_inst38_o0 = inverter1n_inst3_o0 & phasebus_0;
  assign and2n_inst39_o0 = cmpp_eq_inst20_o1 & phasebus_0;
  assign and2n_inst40_o0 = cmpp_eq_inst20_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst1(
                      .enable0(or3n_inst1_o0),
                      .enable1(and2n_inst42_o0),
                      .i0(select_2_1_wn_inst2_o0[11 : 0]),
                      .i1(12'b000000000000),
                      .o0(select_2_1_wn_inst1_o0[11 : 0]));

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst2(
                      .enable0(and2n_inst39_o0),
                      .enable1(and2n_inst40_o0),
                      .i0(addw_inst3_o0[11 : 0]),
                      .i1(sext_inst71_o0[11 : 0]),
                      .o0(select_2_1_wn_inst2_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst71(
                      .i0(1'b0),
                      .o0(sext_inst71_o0[11 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:15  
  sregn_noinitreset #(.width(12))  rr_var_x_stage_3(
                      .clk(clk),
                      .enable(and2n_inst44_o0),
                      .i0(select_2_1_wn_inst1_o0[11 : 0]),
                      .o0(rr_var_x_stage_3_o0[11 : 0]));

  assign and2n_inst41_o0 = or3n_inst2_o0 & and3n_inst0_o0;
  assign inverter1n_inst4_o0 = ~or3n_inst1_o0;
  assign and2n_inst42_o0 = sig_start & inverter1n_inst4_o0;
  assign or3n_inst3_o0 = and2n_inst38_o0 | and2n_inst39_o0 | and2n_inst40_o0;
  assign inverter1n_inst5_o0 = ~and2n_inst43_o0;
  assign and2n_inst43_o0 = and2n_inst38_o0 & or3n_inst3_o0;
  assign and2n_inst44_o0 = and2n_inst41_o0 & inverter1n_inst5_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:15  
  sregn_noinitreset #(.width(12))  rr_var_x_stage_4(
                      .clk(clk),
                      .enable(and2n_inst45_o0),
                      .i0(rr_var_x_stage_3_o0[11 : 0]),
                      .o0(rr_var_x_stage_4_o0[11 : 0]));

  assign and2n_inst45_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:15  
  sregn_noinitreset #(.width(12))  rr_var_x_stage_5(
                      .clk(clk),
                      .enable(and2n_inst46_o0),
                      .i0(rr_var_x_stage_4_o0[11 : 0]),
                      .o0(rr_var_x_stage_5_o0[11 : 0]));

  assign and2n_inst46_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:15  
  sregn_noinitreset #(.width(12))  rr_var_x_stage_6(
                      .clk(clk),
                      .enable(and2n_inst47_o0),
                      .i0(rr_var_x_stage_5_o0[11 : 0]),
                      .o0(rr_var_x_stage_6_o0[11 : 0]));

  assign and2n_inst47_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:15  
  sregn_noinitreset #(.width(12))  rr_var_x_stage_7(
                      .clk(clk),
                      .enable(and2n_inst48_o0),
                      .i0(rr_var_x_stage_6_o0[11 : 0]),
                      .o0(rr_var_x_stage_7_o0[11 : 0]));

  assign and2n_inst48_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:15  
  sregn_noinitreset #(.width(12))  rr_var_x_stage_8(
                      .clk(clk),
                      .enable(and2n_inst49_o0),
                      .i0(rr_var_x_stage_7_o0[11 : 0]),
                      .o0(rr_var_x_stage_8_o0[11 : 0]));

  assign and2n_inst49_o0 = phasebus_0 & and3n_inst0_o0;
  assign or2n_inst9_o0 = and2n_inst50_o0 | and2n_inst51_o0;
  assign or3n_inst4_o0 = and2n_inst51_o0 | sig_start | phasebus_0;
  assign inverter1n_inst6_o0 = ~and2n_inst51_o0;
  assign and2n_inst50_o0 = inverter1n_inst6_o0 & phasebus_0;
  assign and2n_inst51_o0 = rr_func_cmpp_eq_inst12_0_stage_5_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(1))  select_2_1_wn_inst3(
                      .enable0(or2n_inst9_o0),
                      .enable1(and2n_inst53_o0),
                      .i0(datamerge_select_2_1_wn_inst25_o0),
                      .i1(1'b0),
                      .o0(select_2_1_wn_inst3_o0));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst55_o0),
                      .i0(select_2_1_wn_inst3_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_6_o0));

  assign and2n_inst52_o0 = or3n_inst4_o0 & and3n_inst0_o0;
  assign inverter1n_inst7_o0 = ~or2n_inst9_o0;
  assign and2n_inst53_o0 = sig_start & inverter1n_inst7_o0;
  assign or2n_inst11_o0 = and2n_inst50_o0 | and2n_inst51_o0;
  assign nor2n_inst0_o0 = ~(and3n_inst1_o0 | and2n_inst54_o0);
  assign and3n_inst1_o0 = nor2n_inst3_o0 & and2n_inst51_o0 & or2n_inst11_o0;
  assign and2n_inst54_o0 = and2n_inst50_o0 & or2n_inst11_o0;
  assign and2n_inst55_o0 = and2n_inst52_o0 & nor2n_inst0_o0;
  assign or2n_inst12_o0 = and2n_inst58_o0 | and2n_inst57_o0;
  assign or2n_inst13_o0 = or2n_inst12_o0 | phasebus_0;
  assign inverter1n_inst8_o0 = ~or2n_inst12_o0;
  assign and2n_inst56_o0 = inverter1n_inst8_o0 & phasebus_0;
  assign and2n_inst57_o0 = rr_func_cmpp_eq_inst12_stage_6_o0 & phasebus_0;
  assign and2n_inst58_o0 = rr_func_cmpp_eq_inst0_stage_6_o0 & phasebus_0;

  select_3_1_wn #(.dwidth(1))  select_3_1_wn_inst1(
                      .enable0(and2n_inst56_o0),
                      .enable1(and2n_inst57_o0),
                      .enable2(and2n_inst58_o0),
                      .i0(rr_var_dvi_ds_s_hs_stage_6_o0),
                      .i1(datamerge_select_2_1_wn_inst26_o0[0]),
                      .i2(datamerge_select_2_1_wn_inst24_o0[0]),
                      .o0(select_3_1_wn_inst1_o0));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst59_o0),
                      .i0(select_3_1_wn_inst1_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_7_o0));

  assign and2n_inst59_o0 = or2n_inst13_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst60_o0),
                      .i0(rr_var_dvi_ds_s_hs_stage_7_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_8_o0));

  assign and2n_inst60_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst61_o0),
                      .i0(rr_var_dvi_ds_s_hs_stage_8_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_9_o0));

  assign and2n_inst61_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst62_o0),
                      .i0(rr_var_dvi_ds_s_hs_stage_9_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_10_o0));

  assign and2n_inst62_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst63_o0),
                      .i0(rr_var_dvi_ds_s_hs_stage_10_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_11_o0));

  assign and2n_inst63_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_hs_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst64_o0),
                      .i0(rr_var_dvi_ds_s_hs_stage_11_o0),
                      .o0(rr_var_dvi_ds_s_hs_stage_12_o0));

  assign and2n_inst64_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst65_o0 = cmpp_eq_inst12_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst66_o0),
                      .i0(cmpp_eq_inst12_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_4_o0));

  assign and2n_inst66_o0 = and2n_inst65_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst67_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_5_o0));

  assign and2n_inst67_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst68_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_6_o0));

  assign and2n_inst68_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst69_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_7_o0));

  assign and2n_inst69_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst70_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_8_o0));

  assign and2n_inst70_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst71_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_9_o0));

  assign and2n_inst71_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst72_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_10_o0));

  assign and2n_inst72_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst73_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_11_o0));

  assign and2n_inst73_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst74_o0),
                      .i0(rr_func_cmpp_eq_inst12_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst12_stage_12_o0));

  assign and2n_inst74_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst75_o0 = cmpp_eq_inst12_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_0_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst76_o0),
                      .i0(cmpp_eq_inst12_o1),
                      .o0(rr_func_cmpp_eq_inst12_0_stage_4_o0));

  assign and2n_inst76_o0 = and2n_inst75_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:74:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst12_0_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst77_o0),
                      .i0(rr_func_cmpp_eq_inst12_0_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst12_0_stage_5_o0));

  assign and2n_inst77_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst78_o0 = addw_inst4_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:25  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:25  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst4_stage_5(
                      .clk(clk),
                      .enable(and2n_inst79_o0),
                      .i0(addw_inst4_o0[31 : 0]),
                      .o0(rr_func_addw_inst4_stage_5_o0[31 : 0]));

  assign and2n_inst79_o0 = and2n_inst78_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:25  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:25  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst4_stage_6(
                      .clk(clk),
                      .enable(and2n_inst80_o0),
                      .i0(rr_func_addw_inst4_stage_5_o0[31 : 0]),
                      .o0(rr_func_addw_inst4_stage_6_o0[31 : 0]));

  assign and2n_inst80_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst81_o0 = cmpp_eq_inst13_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst82_o0),
                      .i0(cmpp_eq_inst13_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_6_o0));

  assign and2n_inst82_o0 = and2n_inst81_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst83_o0),
                      .i0(rr_func_cmpp_eq_inst13_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_7_o0));

  assign and2n_inst83_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst84_o0),
                      .i0(rr_func_cmpp_eq_inst13_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_8_o0));

  assign and2n_inst84_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst85_o0),
                      .i0(rr_func_cmpp_eq_inst13_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_9_o0));

  assign and2n_inst85_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst86_o0),
                      .i0(rr_func_cmpp_eq_inst13_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_10_o0));

  assign and2n_inst86_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst87_o0),
                      .i0(rr_func_cmpp_eq_inst13_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_11_o0));

  assign and2n_inst87_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst88_o0),
                      .i0(rr_func_cmpp_eq_inst13_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst13_stage_12_o0));

  assign and2n_inst88_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst89_o0 = cmpp_eq_inst13_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_0_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst90_o0),
                      .i0(cmpp_eq_inst13_o1),
                      .o0(rr_func_cmpp_eq_inst13_0_stage_6_o0));

  assign and2n_inst90_o0 = and2n_inst89_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:76:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst13_0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst91_o0),
                      .i0(rr_func_cmpp_eq_inst13_0_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst13_0_stage_7_o0));

  assign and2n_inst91_o0 = phasebus_0 & and3n_inst0_o0;
  assign or3n_inst6_o0 = and2n_inst92_o0 | and2n_inst93_o0 | and2n_inst94_o0;
  assign or3n_inst7_o0 = and2n_inst95_o0 | and2n_inst96_o0 | and2n_inst97_o0;
  assign or2n_inst14_o0 = or3n_inst6_o0 | or3n_inst7_o0;
  assign or3n_inst8_o0 = and2n_inst97_o0 | and2n_inst93_o0 | and2n_inst94_o0;
  assign or2n_inst15_o0 = and2n_inst95_o0 | and2n_inst96_o0;
  assign or2n_inst16_o0 = or3n_inst8_o0 | or2n_inst15_o0;
  assign or3n_inst9_o0 = or2n_inst16_o0 | sig_start | phasebus_0;
  assign inverter1n_inst9_o0 = ~or2n_inst16_o0;
  assign and2n_inst92_o0 = inverter1n_inst9_o0 & phasebus_0;
  assign and2n_inst93_o0 = rr_func_cmpp_eq_inst14_stage_12_o0 & phasebus_0;
  assign and2n_inst94_o0 = rr_func_cmpp_eq_inst14_0_stage_12_o0 & phasebus_0;
  assign and2n_inst95_o0 = rr_func_cmpp_eq_inst0_stage_12_o0 & phasebus_0;
  assign and2n_inst96_o0 = rr_func_cmpp_eq_inst12_stage_12_o0 & phasebus_0;
  assign and2n_inst97_o0 = rr_func_cmpp_eq_inst13_stage_12_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst4(
                      .enable0(or2n_inst14_o0),
                      .enable1(and2n_inst99_o0),
                      .i0(select_2_1_wn_inst5_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst4_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst5(
                      .enable0(and2n_inst93_o0),
                      .enable1(and2n_inst97_o0),
                      .i0(sext_inst72_o0[1 : 0]),
                      .i1(sext_inst19_o0[1 : 0]),
                      .o0(select_2_1_wn_inst5_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst72(
                      .i0(1'b0),
                      .o0(sext_inst72_o0[1 : 0]));

  assign or3n_inst10_o0 = and2n_inst94_o0 | and2n_inst95_o0 | and2n_inst96_o0;
  assign or2n_inst19_o0 = or3n_inst10_o0 | and2n_inst92_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:68:7  
  sregn_noinitreset #(.width(2))  rr_var_hactive_stage_13(
                      .clk(clk),
                      .enable(and2n_inst101_o0),
                      .i0(select_2_1_wn_inst4_o0[1 : 0]),
                      .o0(rr_var_hactive_stage_13_o0[1 : 0]));

  assign and2n_inst98_o0 = or3n_inst9_o0 & and3n_inst0_o0;
  assign inverter1n_inst10_o0 = ~or2n_inst14_o0;
  assign and2n_inst99_o0 = sig_start & inverter1n_inst10_o0;
  assign or3n_inst11_o0 = and2n_inst92_o0 | and2n_inst93_o0 | and2n_inst94_o0;
  assign or3n_inst12_o0 = and2n_inst95_o0 | and2n_inst96_o0 | and2n_inst97_o0;
  assign or2n_inst20_o0 = or3n_inst11_o0 | or3n_inst12_o0;
  assign inverter1n_inst11_o0 = ~and2n_inst100_o0;
  assign and2n_inst100_o0 = or2n_inst19_o0 & or2n_inst20_o0;
  assign and2n_inst101_o0 = and2n_inst98_o0 & inverter1n_inst11_o0;
  assign and2n_inst102_o0 = addw_inst5_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:35  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst5_stage_7(
                      .clk(clk),
                      .enable(and2n_inst103_o0),
                      .i0(addw_inst5_o0[31 : 0]),
                      .o0(rr_func_addw_inst5_stage_7_o0[31 : 0]));

  assign and2n_inst103_o0 = and2n_inst102_o0 & and3n_inst0_o0;
  assign and2n_inst104_o0 = cmpp_eq_inst14_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst105_o0),
                      .i0(cmpp_eq_inst14_o0),
                      .o0(rr_func_cmpp_eq_inst14_stage_8_o0));

  assign and2n_inst105_o0 = and2n_inst104_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst106_o0),
                      .i0(rr_func_cmpp_eq_inst14_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst14_stage_9_o0));

  assign and2n_inst106_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst107_o0),
                      .i0(rr_func_cmpp_eq_inst14_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst14_stage_10_o0));

  assign and2n_inst107_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst108_o0),
                      .i0(rr_func_cmpp_eq_inst14_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst14_stage_11_o0));

  assign and2n_inst108_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst109_o0),
                      .i0(rr_func_cmpp_eq_inst14_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst14_stage_12_o0));

  assign and2n_inst109_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst110_o0 = cmpp_eq_inst14_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_0_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst111_o0),
                      .i0(cmpp_eq_inst14_o1),
                      .o0(rr_func_cmpp_eq_inst14_0_stage_8_o0));

  assign and2n_inst111_o0 = and2n_inst110_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_0_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst112_o0),
                      .i0(rr_func_cmpp_eq_inst14_0_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst14_0_stage_9_o0));

  assign and2n_inst112_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst113_o0),
                      .i0(rr_func_cmpp_eq_inst14_0_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst14_0_stage_10_o0));

  assign and2n_inst113_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst114_o0),
                      .i0(rr_func_cmpp_eq_inst14_0_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst14_0_stage_11_o0));

  assign and2n_inst114_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:78:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst14_0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst115_o0),
                      .i0(rr_func_cmpp_eq_inst14_0_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst14_0_stage_12_o0));

  assign and2n_inst115_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst116_o0 = cmpp_eq_inst1_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst117_o0),
                      .i0(cmpp_eq_inst1_o0),
                      .o0(rr_func_cmpp_eq_inst1_stage_7_o0));

  assign and2n_inst117_o0 = and2n_inst116_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst118_o0),
                      .i0(rr_func_cmpp_eq_inst1_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst1_stage_8_o0));

  assign and2n_inst118_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst119_o0),
                      .i0(rr_func_cmpp_eq_inst1_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst1_stage_9_o0));

  assign and2n_inst119_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst120_o0),
                      .i0(rr_func_cmpp_eq_inst1_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst1_stage_10_o0));

  assign and2n_inst120_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst121_o0),
                      .i0(rr_func_cmpp_eq_inst1_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst1_stage_11_o0));

  assign and2n_inst121_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst122_o0),
                      .i0(rr_func_cmpp_eq_inst1_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst1_stage_12_o0));

  assign and2n_inst122_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst123_o0 = cmpp_eq_inst1_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:82:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst1_0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst124_o0),
                      .i0(cmpp_eq_inst1_o1),
                      .o0(rr_func_cmpp_eq_inst1_0_stage_7_o0));

  assign and2n_inst124_o0 = and2n_inst123_o0 & and3n_inst0_o0;
  assign or3n_inst13_o0 = and2n_inst125_o0 | and2n_inst126_o0 | and2n_inst127_o0;
  assign or2n_inst21_o0 = or3n_inst13_o0 | and2n_inst128_o0;
  assign or3n_inst14_o0 = and2n_inst128_o0 | and2n_inst126_o0 | and2n_inst127_o0;
  assign or3n_inst15_o0 = or3n_inst14_o0 | sig_start | phasebus_0;
  assign inverter1n_inst12_o0 = ~or3n_inst14_o0;
  assign and2n_inst125_o0 = inverter1n_inst12_o0 & phasebus_0;
  assign and2n_inst126_o0 = cmpp_eq_inst21_o1 & phasebus_0;
  assign and2n_inst127_o0 = rr_func_cmpp_eq_inst20_0_stage_6_o0 & phasebus_0;
  assign and2n_inst128_o0 = cmpp_eq_inst21_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst6(
                      .enable0(or2n_inst21_o0),
                      .enable1(and2n_inst130_o0),
                      .i0(select_2_1_wn_inst7_o0[11 : 0]),
                      .i1(12'b000000000000),
                      .o0(select_2_1_wn_inst6_o0[11 : 0]));

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst7(
                      .enable0(and2n_inst126_o0),
                      .enable1(and2n_inst128_o0),
                      .i0(addw_inst1_o0[11 : 0]),
                      .i1(sext_inst73_o0[11 : 0]),
                      .o0(select_2_1_wn_inst7_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst73(
                      .i0(1'b0),
                      .o0(sext_inst73_o0[11 : 0]));

  assign or2n_inst24_o0 = and2n_inst127_o0 | and2n_inst125_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:22  
  sregn_noinitreset #(.width(12))  rr_var_y_stage_7(
                      .clk(clk),
                      .enable(and2n_inst132_o0),
                      .i0(select_2_1_wn_inst6_o0[11 : 0]),
                      .o0(rr_var_y_stage_7_o0[11 : 0]));

  assign and2n_inst129_o0 = or3n_inst15_o0 & and3n_inst0_o0;
  assign inverter1n_inst13_o0 = ~or2n_inst21_o0;
  assign and2n_inst130_o0 = sig_start & inverter1n_inst13_o0;
  assign or3n_inst16_o0 = and2n_inst125_o0 | and2n_inst126_o0 | and2n_inst127_o0;
  assign or2n_inst25_o0 = or3n_inst16_o0 | and2n_inst128_o0;
  assign inverter1n_inst14_o0 = ~and2n_inst131_o0;
  assign and2n_inst131_o0 = or2n_inst24_o0 & or2n_inst25_o0;
  assign and2n_inst132_o0 = and2n_inst129_o0 & inverter1n_inst14_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:22  
  sregn_noinitreset #(.width(12))  rr_var_y_stage_8(
                      .clk(clk),
                      .enable(and2n_inst133_o0),
                      .i0(rr_var_y_stage_7_o0[11 : 0]),
                      .o0(rr_var_y_stage_8_o0[11 : 0]));

  assign and2n_inst133_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:22  
  sregn_noinitreset #(.width(12))  rr_var_y_stage_9(
                      .clk(clk),
                      .enable(and2n_inst134_o0),
                      .i0(rr_var_y_stage_8_o0[11 : 0]),
                      .o0(rr_var_y_stage_9_o0[11 : 0]));

  assign and2n_inst134_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:22  
  sregn_noinitreset #(.width(12))  rr_var_y_stage_10(
                      .clk(clk),
                      .enable(and2n_inst135_o0),
                      .i0(rr_var_y_stage_9_o0[11 : 0]),
                      .o0(rr_var_y_stage_10_o0[11 : 0]));

  assign and2n_inst135_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:22  
  sregn_noinitreset #(.width(12))  rr_var_y_stage_11(
                      .clk(clk),
                      .enable(and2n_inst136_o0),
                      .i0(rr_var_y_stage_10_o0[11 : 0]),
                      .o0(rr_var_y_stage_11_o0[11 : 0]));

  assign and2n_inst136_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:62:22  
  sregn_noinitreset #(.width(12))  rr_var_y_stage_12(
                      .clk(clk),
                      .enable(and2n_inst137_o0),
                      .i0(rr_var_y_stage_11_o0[11 : 0]),
                      .o0(rr_var_y_stage_12_o0[11 : 0]));

  assign and2n_inst137_o0 = phasebus_0 & and3n_inst0_o0;
  assign or2n_inst26_o0 = and2n_inst138_o0 | and2n_inst139_o0;
  assign or3n_inst17_o0 = and2n_inst139_o0 | sig_start | phasebus_0;
  assign inverter1n_inst15_o0 = ~and2n_inst139_o0;
  assign and2n_inst138_o0 = inverter1n_inst15_o0 & phasebus_0;
  assign and2n_inst139_o0 = rr_func_cmpp_eq_inst15_0_stage_11_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(1))  select_2_1_wn_inst8(
                      .enable0(or2n_inst26_o0),
                      .enable1(and2n_inst141_o0),
                      .i0(datamerge_select_2_1_wn_inst28_o0),
                      .i1(1'b0),
                      .o0(select_2_1_wn_inst8_o0));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:70:18  
  sregn_noinit #(.width(1))  rr_var_dvi_ds_s_vs_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst143_o0),
                      .i0(select_2_1_wn_inst8_o0),
                      .o0(rr_var_dvi_ds_s_vs_stage_12_o0));

  assign and2n_inst140_o0 = or3n_inst17_o0 & and3n_inst0_o0;
  assign inverter1n_inst16_o0 = ~or2n_inst26_o0;
  assign and2n_inst141_o0 = sig_start & inverter1n_inst16_o0;
  assign or2n_inst28_o0 = and2n_inst138_o0 | and2n_inst139_o0;
  assign nor2n_inst1_o0 = ~(and3n_inst2_o0 | and2n_inst142_o0);
  assign and3n_inst2_o0 = nor2n_inst5_o0 & and2n_inst139_o0 & or2n_inst28_o0;
  assign and2n_inst142_o0 = and2n_inst138_o0 & or2n_inst28_o0;
  assign and2n_inst143_o0 = and2n_inst140_o0 & nor2n_inst1_o0;
  assign and2n_inst144_o0 = cmpp_eq_inst15_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst145_o0),
                      .i0(cmpp_eq_inst15_o0),
                      .o0(rr_func_cmpp_eq_inst15_stage_8_o0));

  assign and2n_inst145_o0 = and2n_inst144_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst146_o0),
                      .i0(rr_func_cmpp_eq_inst15_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst15_stage_9_o0));

  assign and2n_inst146_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst147_o0),
                      .i0(rr_func_cmpp_eq_inst15_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst15_stage_10_o0));

  assign and2n_inst147_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst148_o0),
                      .i0(rr_func_cmpp_eq_inst15_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst15_stage_11_o0));

  assign and2n_inst148_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst149_o0),
                      .i0(rr_func_cmpp_eq_inst15_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst15_stage_12_o0));

  assign and2n_inst149_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst150_o0 = cmpp_eq_inst15_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_0_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst151_o0),
                      .i0(cmpp_eq_inst15_o1),
                      .o0(rr_func_cmpp_eq_inst15_0_stage_8_o0));

  assign and2n_inst151_o0 = and2n_inst150_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_0_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst152_o0),
                      .i0(rr_func_cmpp_eq_inst15_0_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst15_0_stage_9_o0));

  assign and2n_inst152_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst153_o0),
                      .i0(rr_func_cmpp_eq_inst15_0_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst15_0_stage_10_o0));

  assign and2n_inst153_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:84:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst15_0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst154_o0),
                      .i0(rr_func_cmpp_eq_inst15_0_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst15_0_stage_11_o0));

  assign and2n_inst154_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst155_o0 = addw_inst6_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:25  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:25  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst6_stage_9(
                      .clk(clk),
                      .enable(and2n_inst156_o0),
                      .i0(addw_inst6_o0[31 : 0]),
                      .o0(rr_func_addw_inst6_stage_9_o0[31 : 0]));

  assign and2n_inst156_o0 = and2n_inst155_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:25  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:25  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst6_stage_10(
                      .clk(clk),
                      .enable(and2n_inst157_o0),
                      .i0(rr_func_addw_inst6_stage_9_o0[31 : 0]),
                      .o0(rr_func_addw_inst6_stage_10_o0[31 : 0]));

  assign and2n_inst157_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst158_o0 = cmpp_eq_inst16_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst16_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst159_o0),
                      .i0(cmpp_eq_inst16_o0),
                      .o0(rr_func_cmpp_eq_inst16_stage_10_o0));

  assign and2n_inst159_o0 = and2n_inst158_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst16_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst160_o0),
                      .i0(rr_func_cmpp_eq_inst16_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst16_stage_11_o0));

  assign and2n_inst160_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst16_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst161_o0),
                      .i0(rr_func_cmpp_eq_inst16_stage_11_o0),
                      .o0(rr_func_cmpp_eq_inst16_stage_12_o0));

  assign and2n_inst161_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst162_o0 = cmpp_eq_inst16_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst16_0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst163_o0),
                      .i0(cmpp_eq_inst16_o1),
                      .o0(rr_func_cmpp_eq_inst16_0_stage_10_o0));

  assign and2n_inst163_o0 = and2n_inst162_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:86:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst16_0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst164_o0),
                      .i0(rr_func_cmpp_eq_inst16_0_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst16_0_stage_11_o0));

  assign and2n_inst164_o0 = phasebus_0 & and3n_inst0_o0;
  assign or3n_inst18_o0 = and2n_inst165_o0 | and2n_inst166_o0 | and2n_inst167_o0;
  assign or3n_inst19_o0 = and2n_inst168_o0 | and2n_inst169_o0 | and2n_inst170_o0;
  assign or2n_inst29_o0 = or3n_inst18_o0 | or3n_inst19_o0;
  assign or3n_inst20_o0 = and2n_inst170_o0 | and2n_inst166_o0 | and2n_inst167_o0;
  assign or2n_inst30_o0 = and2n_inst168_o0 | and2n_inst169_o0;
  assign or2n_inst31_o0 = or3n_inst20_o0 | or2n_inst30_o0;
  assign or3n_inst21_o0 = or2n_inst31_o0 | sig_start | phasebus_0;
  assign inverter1n_inst17_o0 = ~or2n_inst31_o0;
  assign and2n_inst165_o0 = inverter1n_inst17_o0 & phasebus_0;
  assign and2n_inst166_o0 = rr_func_cmpp_eq_inst17_stage_12_o0 & phasebus_0;
  assign and2n_inst167_o0 = rr_func_cmpp_eq_inst17_0_stage_12_o0 & phasebus_0;
  assign and2n_inst168_o0 = rr_func_cmpp_eq_inst1_stage_12_o0 & phasebus_0;
  assign and2n_inst169_o0 = rr_func_cmpp_eq_inst15_stage_12_o0 & phasebus_0;
  assign and2n_inst170_o0 = rr_func_cmpp_eq_inst16_stage_12_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst9(
                      .enable0(or2n_inst29_o0),
                      .enable1(and2n_inst172_o0),
                      .i0(select_2_1_wn_inst10_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst9_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst10(
                      .enable0(and2n_inst166_o0),
                      .enable1(and2n_inst170_o0),
                      .i0(sext_inst74_o0[1 : 0]),
                      .i1(sext_inst23_o0[1 : 0]),
                      .o0(select_2_1_wn_inst10_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst74(
                      .i0(1'b0),
                      .o0(sext_inst74_o0[1 : 0]));

  assign or3n_inst22_o0 = and2n_inst167_o0 | and2n_inst168_o0 | and2n_inst169_o0;
  assign or2n_inst34_o0 = or3n_inst22_o0 | and2n_inst165_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:68:19  
  sregn_noinitreset #(.width(2))  rr_var_vactive_stage_13(
                      .clk(clk),
                      .enable(and2n_inst174_o0),
                      .i0(select_2_1_wn_inst9_o0[1 : 0]),
                      .o0(rr_var_vactive_stage_13_o0[1 : 0]));

  assign and2n_inst171_o0 = or3n_inst21_o0 & and3n_inst0_o0;
  assign inverter1n_inst18_o0 = ~or2n_inst29_o0;
  assign and2n_inst172_o0 = sig_start & inverter1n_inst18_o0;
  assign or3n_inst23_o0 = and2n_inst165_o0 | and2n_inst166_o0 | and2n_inst167_o0;
  assign or3n_inst24_o0 = and2n_inst168_o0 | and2n_inst169_o0 | and2n_inst170_o0;
  assign or2n_inst35_o0 = or3n_inst23_o0 | or3n_inst24_o0;
  assign inverter1n_inst19_o0 = ~and2n_inst173_o0;
  assign and2n_inst173_o0 = or2n_inst34_o0 & or2n_inst35_o0;
  assign and2n_inst174_o0 = and2n_inst171_o0 & inverter1n_inst19_o0;
  assign and2n_inst175_o0 = addw_inst7_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:35  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst7_stage_11(
                      .clk(clk),
                      .enable(and2n_inst176_o0),
                      .i0(addw_inst7_o0[31 : 0]),
                      .o0(rr_func_addw_inst7_stage_11_o0[31 : 0]));

  assign and2n_inst176_o0 = and2n_inst175_o0 & and3n_inst0_o0;
  assign and2n_inst177_o0 = cmpp_eq_inst17_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst17_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst178_o0),
                      .i0(cmpp_eq_inst17_o0),
                      .o0(rr_func_cmpp_eq_inst17_stage_12_o0));

  assign and2n_inst178_o0 = and2n_inst177_o0 & and3n_inst0_o0;
  assign and2n_inst179_o0 = cmpp_eq_inst17_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:88:15  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst17_0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst180_o0),
                      .i0(cmpp_eq_inst17_o1),
                      .o0(rr_func_cmpp_eq_inst17_0_stage_12_o0));

  assign and2n_inst180_o0 = and2n_inst179_o0 & and3n_inst0_o0;
  assign and2n_inst181_o0 = addw_inst8_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:18  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:28  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst8_stage_0(
                      .clk(clk),
                      .enable(and2n_inst182_o0),
                      .i0(addw_inst8_o0[31 : 0]),
                      .o0(rr_func_addw_inst8_stage_0_o0[31 : 0]));

  assign and2n_inst182_o0 = and2n_inst181_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:18  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:28  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst8_stage_1(
                      .clk(clk),
                      .enable(and2n_inst183_o0),
                      .i0(rr_func_addw_inst8_stage_0_o0[31 : 0]),
                      .o0(rr_func_addw_inst8_stage_1_o0[31 : 0]));

  assign and2n_inst183_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:18  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:28  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst8_stage_2(
                      .clk(clk),
                      .enable(and2n_inst184_o0),
                      .i0(rr_func_addw_inst8_stage_1_o0[31 : 0]),
                      .o0(rr_func_addw_inst8_stage_2_o0[31 : 0]));

  assign and2n_inst184_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst185_o0 = cmpp_eq_inst18_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst186_o0),
                      .i0(cmpp_eq_inst18_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_3_o0));

  assign and2n_inst186_o0 = and2n_inst185_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst187_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_3_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_4_o0));

  assign and2n_inst187_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst188_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_5_o0));

  assign and2n_inst188_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst189_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_6_o0));

  assign and2n_inst189_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst190_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_7_o0));

  assign and2n_inst190_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst191_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_8_o0));

  assign and2n_inst191_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst192_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_9_o0));

  assign and2n_inst192_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst193_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_10_o0));

  assign and2n_inst193_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst194_o0),
                      .i0(rr_func_cmpp_eq_inst18_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst18_stage_11_o0));

  assign and2n_inst194_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst195_o0 = cmpp_eq_inst18_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:92:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst18_0_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst196_o0),
                      .i0(cmpp_eq_inst18_o1),
                      .o0(rr_func_cmpp_eq_inst18_0_stage_3_o0));

  assign and2n_inst196_o0 = and2n_inst195_o0 & and3n_inst0_o0;
  assign or3n_inst25_o0 = and2n_inst197_o0 | and2n_inst198_o0 | and2n_inst199_o0;
  assign or2n_inst36_o0 = and2n_inst199_o0 | and2n_inst198_o0;
  assign or3n_inst26_o0 = or2n_inst36_o0 | sig_start | phasebus_0;
  assign inverter1n_inst20_o0 = ~or2n_inst36_o0;
  assign and2n_inst197_o0 = inverter1n_inst20_o0 & phasebus_0;
  assign and2n_inst198_o0 = cmpp_eq_inst22_o1 & phasebus_0;
  assign and2n_inst199_o0 = cmpp_eq_inst22_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst11(
                      .enable0(or3n_inst25_o0),
                      .enable1(and2n_inst201_o0),
                      .i0(select_2_1_wn_inst12_o0[11 : 0]),
                      .i1(12'b000000000000),
                      .o0(select_2_1_wn_inst11_o0[11 : 0]));

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst12(
                      .enable0(and2n_inst198_o0),
                      .enable1(and2n_inst199_o0),
                      .i0(addw_inst0_o0[11 : 0]),
                      .i1(sext_inst75_o0[11 : 0]),
                      .o0(select_2_1_wn_inst12_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst75(
                      .i0(1'b0),
                      .o0(sext_inst75_o0[11 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:65:15  
  sregn_noinitreset #(.width(12))  rr_var_xa_stage_4(
                      .clk(clk),
                      .enable(and2n_inst203_o0),
                      .i0(select_2_1_wn_inst11_o0[11 : 0]),
                      .o0(rr_var_xa_stage_4_o0[11 : 0]));

  assign and2n_inst200_o0 = or3n_inst26_o0 & and3n_inst0_o0;
  assign inverter1n_inst21_o0 = ~or3n_inst25_o0;
  assign and2n_inst201_o0 = sig_start & inverter1n_inst21_o0;
  assign or3n_inst27_o0 = and2n_inst197_o0 | and2n_inst198_o0 | and2n_inst199_o0;
  assign inverter1n_inst22_o0 = ~and2n_inst202_o0;
  assign and2n_inst202_o0 = and2n_inst197_o0 & or3n_inst27_o0;
  assign and2n_inst203_o0 = and2n_inst200_o0 & inverter1n_inst22_o0;
  assign or3n_inst28_o0 = and2n_inst204_o0 | and2n_inst205_o0 | and2n_inst206_o0;
  assign or2n_inst39_o0 = or3n_inst28_o0 | and2n_inst207_o0;
  assign or3n_inst29_o0 = and2n_inst207_o0 | and2n_inst205_o0 | and2n_inst206_o0;
  assign or3n_inst30_o0 = or3n_inst29_o0 | sig_start | phasebus_0;
  assign inverter1n_inst23_o0 = ~or3n_inst29_o0;
  assign and2n_inst204_o0 = inverter1n_inst23_o0 & phasebus_0;
  assign and2n_inst205_o0 = rr_func_cmpp_eq_inst22_stage_11_o0 & phasebus_0;
  assign and2n_inst206_o0 = rr_func_cmpp_eq_inst22_0_stage_11_o0 & phasebus_0;
  assign and2n_inst207_o0 = rr_func_cmpp_eq_inst18_stage_11_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst13(
                      .enable0(or2n_inst39_o0),
                      .enable1(and2n_inst209_o0),
                      .i0(select_2_1_wn_inst14_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst13_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst14(
                      .enable0(and2n_inst205_o0),
                      .enable1(and2n_inst207_o0),
                      .i0(rr_func_moveii_inst40_stage_11_o0[1 : 0]),
                      .i1(sext_inst24_o0[1 : 0]),
                      .o0(select_2_1_wn_inst14_o0[1 : 0]));

  assign or2n_inst42_o0 = and2n_inst206_o0 | and2n_inst204_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:69:66  
  sregn_noinitreset #(.width(2))  rr_var_bactive_stage_12(
                      .clk(clk),
                      .enable(and2n_inst211_o0),
                      .i0(select_2_1_wn_inst13_o0[1 : 0]),
                      .o0(rr_var_bactive_stage_12_o0[1 : 0]));

  assign and2n_inst208_o0 = or3n_inst30_o0 & and3n_inst0_o0;
  assign inverter1n_inst24_o0 = ~or2n_inst39_o0;
  assign and2n_inst209_o0 = sig_start & inverter1n_inst24_o0;
  assign or3n_inst31_o0 = and2n_inst204_o0 | and2n_inst205_o0 | and2n_inst206_o0;
  assign or2n_inst43_o0 = or3n_inst31_o0 | and2n_inst207_o0;
  assign inverter1n_inst25_o0 = ~and2n_inst210_o0;
  assign and2n_inst210_o0 = or2n_inst42_o0 & or2n_inst43_o0;
  assign and2n_inst211_o0 = and2n_inst208_o0 & inverter1n_inst25_o0;
  assign or3n_inst32_o0 = and2n_inst212_o0 | and2n_inst213_o0 | and2n_inst214_o0;
  assign or2n_inst44_o0 = and2n_inst215_o0 | and2n_inst216_o0;
  assign or2n_inst45_o0 = or3n_inst32_o0 | or2n_inst44_o0;
  assign or3n_inst33_o0 = and2n_inst216_o0 | and2n_inst213_o0 | and2n_inst214_o0;
  assign or2n_inst46_o0 = or3n_inst33_o0 | and2n_inst215_o0;
  assign or3n_inst34_o0 = or2n_inst46_o0 | sig_start | phasebus_0;
  assign inverter1n_inst26_o0 = ~or2n_inst46_o0;
  assign and2n_inst212_o0 = inverter1n_inst26_o0 & phasebus_0;
  assign and2n_inst213_o0 = cmpp_eq_inst6_o0 & phasebus_0;
  assign and2n_inst214_o0 = rr_func_cmpp_eq_inst22_0_stage_11_o0 & phasebus_0;
  assign and2n_inst215_o0 = cmpp_eq_inst6_o1 & phasebus_0;
  assign and2n_inst216_o0 = rr_func_cmpp_eq_inst18_stage_11_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst15(
                      .enable0(or2n_inst45_o0),
                      .enable1(and2n_inst218_o0),
                      .i0(select_2_1_wn_inst16_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst15_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst16(
                      .enable0(and2n_inst213_o0),
                      .enable1(and2n_inst216_o0),
                      .i0(cmpr_eq_inst2_o0[1 : 0]),
                      .i1(sext_inst25_o0[1 : 0]),
                      .o0(select_2_1_wn_inst16_o0[1 : 0]));

  assign or3n_inst35_o0 = and2n_inst214_o0 | and2n_inst215_o0 | and2n_inst212_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:69:53  
  sregn_noinitreset #(.width(2))  rr_var_gactive_stage_12(
                      .clk(clk),
                      .enable(and2n_inst220_o0),
                      .i0(select_2_1_wn_inst15_o0[1 : 0]),
                      .o0(rr_var_gactive_stage_12_o0[1 : 0]));

  assign and2n_inst217_o0 = or3n_inst34_o0 & and3n_inst0_o0;
  assign inverter1n_inst27_o0 = ~or2n_inst45_o0;
  assign and2n_inst218_o0 = sig_start & inverter1n_inst27_o0;
  assign or3n_inst36_o0 = and2n_inst212_o0 | and2n_inst213_o0 | and2n_inst214_o0;
  assign or2n_inst49_o0 = and2n_inst215_o0 | and2n_inst216_o0;
  assign or2n_inst50_o0 = or3n_inst36_o0 | or2n_inst49_o0;
  assign inverter1n_inst28_o0 = ~and2n_inst219_o0;
  assign and2n_inst219_o0 = or3n_inst35_o0 & or2n_inst50_o0;
  assign and2n_inst220_o0 = and2n_inst217_o0 & inverter1n_inst28_o0;
  assign or3n_inst37_o0 = and2n_inst221_o0 | and2n_inst222_o0 | and2n_inst223_o0;
  assign or2n_inst51_o0 = and2n_inst224_o0 | and2n_inst225_o0;
  assign or2n_inst52_o0 = or3n_inst37_o0 | or2n_inst51_o0;
  assign or3n_inst38_o0 = and2n_inst225_o0 | and2n_inst222_o0 | and2n_inst223_o0;
  assign or2n_inst53_o0 = or3n_inst38_o0 | and2n_inst224_o0;
  assign or3n_inst39_o0 = or2n_inst53_o0 | sig_start | phasebus_0;
  assign inverter1n_inst29_o0 = ~or2n_inst53_o0;
  assign and2n_inst221_o0 = inverter1n_inst29_o0 & phasebus_0;
  assign and2n_inst222_o0 = cmpp_eq_inst7_o0 & phasebus_0;
  assign and2n_inst223_o0 = rr_func_cmpp_eq_inst22_0_stage_11_o0 & phasebus_0;
  assign and2n_inst224_o0 = cmpp_eq_inst7_o1 & phasebus_0;
  assign and2n_inst225_o0 = rr_func_cmpp_eq_inst18_stage_11_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst17(
                      .enable0(or2n_inst52_o0),
                      .enable1(and2n_inst227_o0),
                      .i0(select_2_1_wn_inst18_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst17_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst18(
                      .enable0(and2n_inst222_o0),
                      .enable1(and2n_inst225_o0),
                      .i0(cmpr_eq_inst3_o0[1 : 0]),
                      .i1(sext_inst26_o0[1 : 0]),
                      .o0(select_2_1_wn_inst18_o0[1 : 0]));

  assign or3n_inst40_o0 = and2n_inst223_o0 | and2n_inst224_o0 | and2n_inst221_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:69:40  
  sregn_noinitreset #(.width(2))  rr_var_ractive_stage_12(
                      .clk(clk),
                      .enable(and2n_inst229_o0),
                      .i0(select_2_1_wn_inst17_o0[1 : 0]),
                      .o0(rr_var_ractive_stage_12_o0[1 : 0]));

  assign and2n_inst226_o0 = or3n_inst39_o0 & and3n_inst0_o0;
  assign inverter1n_inst30_o0 = ~or2n_inst52_o0;
  assign and2n_inst227_o0 = sig_start & inverter1n_inst30_o0;
  assign or3n_inst41_o0 = and2n_inst221_o0 | and2n_inst222_o0 | and2n_inst223_o0;
  assign or2n_inst56_o0 = and2n_inst224_o0 | and2n_inst225_o0;
  assign or2n_inst57_o0 = or3n_inst41_o0 | or2n_inst56_o0;
  assign inverter1n_inst31_o0 = ~and2n_inst228_o0;
  assign and2n_inst228_o0 = or3n_inst40_o0 & or2n_inst57_o0;
  assign and2n_inst229_o0 = and2n_inst226_o0 & inverter1n_inst31_o0;
  assign and2n_inst230_o0 = cmpp_eq_inst22_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst231_o0),
                      .i0(cmpp_eq_inst22_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_4_o0));

  assign and2n_inst231_o0 = and2n_inst230_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst232_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_5_o0));

  assign and2n_inst232_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst233_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_6_o0));

  assign and2n_inst233_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst234_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_7_o0));

  assign and2n_inst234_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst235_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_8_o0));

  assign and2n_inst235_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst236_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_9_o0));

  assign and2n_inst236_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst237_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_10_o0));

  assign and2n_inst237_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst238_o0),
                      .i0(rr_func_cmpp_eq_inst22_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst22_stage_11_o0));

  assign and2n_inst238_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst239_o0 = cmpp_eq_inst22_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst240_o0),
                      .i0(cmpp_eq_inst22_o1),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_4_o0));

  assign and2n_inst240_o0 = and2n_inst239_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst241_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_5_o0));

  assign and2n_inst241_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst242_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_6_o0));

  assign and2n_inst242_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst243_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_7_o0));

  assign and2n_inst243_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst244_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_8_o0));

  assign and2n_inst244_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst245_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_9_o0));

  assign and2n_inst245_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst246_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_10_o0));

  assign and2n_inst246_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:97:16  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst22_0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst247_o0),
                      .i0(rr_func_cmpp_eq_inst22_0_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst22_0_stage_11_o0));

  assign and2n_inst247_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst248_o0 = cmpp_neq_inst0_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:7  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst249_o0),
                      .i0(cmpp_neq_inst0_o0),
                      .o0(rr_func_cmpp_neq_inst0_stage_11_o0));

  assign and2n_inst249_o0 = and2n_inst248_o0 & and3n_inst0_o0;
  assign and2n_inst250_o0 = rr_func_cmpp_eq_inst22_stage_10_o0 & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:7  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:104:14  
  sregn_noinitreset #(.width(2))  rr_func_moveii_inst40_stage_11(
                      .clk(clk),
                      .enable(and2n_inst251_o0),
                      .i0(cmpr_eq_inst0_o0[1 : 0]),
                      .o0(rr_func_moveii_inst40_stage_11_o0[1 : 0]));

  assign and2n_inst251_o0 = and2n_inst250_o0 & and3n_inst0_o0;
  assign and2n_inst252_o0 = cmpp_neq_inst0_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:98:7  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst0_0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst253_o0),
                      .i0(cmpp_neq_inst0_o1),
                      .o0(rr_func_cmpp_neq_inst0_0_stage_11_o0));

  assign and2n_inst253_o0 = and2n_inst252_o0 & and3n_inst0_o0;
  assign and2n_inst254_o0 = addw_inst9_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:18  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:29  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst9_stage_4(
                      .clk(clk),
                      .enable(and2n_inst255_o0),
                      .i0(addw_inst9_o0[31 : 0]),
                      .o0(rr_func_addw_inst9_stage_4_o0[31 : 0]));

  assign and2n_inst255_o0 = and2n_inst254_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:18  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:29  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst9_stage_5(
                      .clk(clk),
                      .enable(and2n_inst256_o0),
                      .i0(rr_func_addw_inst9_stage_4_o0[31 : 0]),
                      .o0(rr_func_addw_inst9_stage_5_o0[31 : 0]));

  assign and2n_inst256_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:18  dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:29  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst9_stage_6(
                      .clk(clk),
                      .enable(and2n_inst257_o0),
                      .i0(rr_func_addw_inst9_stage_5_o0[31 : 0]),
                      .o0(rr_func_addw_inst9_stage_6_o0[31 : 0]));

  assign and2n_inst257_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst258_o0 = cmpp_eq_inst19_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst19_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst259_o0),
                      .i0(cmpp_eq_inst19_o0),
                      .o0(rr_func_cmpp_eq_inst19_stage_7_o0));

  assign and2n_inst259_o0 = and2n_inst258_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst19_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst260_o0),
                      .i0(rr_func_cmpp_eq_inst19_stage_7_o0),
                      .o0(rr_func_cmpp_eq_inst19_stage_8_o0));

  assign and2n_inst260_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst19_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst261_o0),
                      .i0(rr_func_cmpp_eq_inst19_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst19_stage_9_o0));

  assign and2n_inst261_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst19_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst262_o0),
                      .i0(rr_func_cmpp_eq_inst19_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst19_stage_10_o0));

  assign and2n_inst262_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst19_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst263_o0),
                      .i0(rr_func_cmpp_eq_inst19_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst19_stage_11_o0));

  assign and2n_inst263_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst264_o0 = cmpp_eq_inst19_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:110:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst19_0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst265_o0),
                      .i0(cmpp_eq_inst19_o1),
                      .o0(rr_func_cmpp_eq_inst19_0_stage_7_o0));

  assign and2n_inst265_o0 = and2n_inst264_o0 & and3n_inst0_o0;
  assign or3n_inst42_o0 = and2n_inst266_o0 | and2n_inst267_o0 | and2n_inst268_o0;
  assign or2n_inst58_o0 = and2n_inst269_o0 | and2n_inst270_o0;
  assign or2n_inst59_o0 = or3n_inst42_o0 | or2n_inst58_o0;
  assign or3n_inst43_o0 = and2n_inst270_o0 | and2n_inst267_o0 | and2n_inst268_o0;
  assign or2n_inst60_o0 = or3n_inst43_o0 | and2n_inst269_o0;
  assign or3n_inst44_o0 = or2n_inst60_o0 | sig_start | phasebus_0;
  assign inverter1n_inst32_o0 = ~or2n_inst60_o0;
  assign and2n_inst266_o0 = inverter1n_inst32_o0 & phasebus_0;
  assign and2n_inst267_o0 = rr_func_cmpp_eq_inst24_stage_10_o0 & phasebus_0;
  assign and2n_inst268_o0 = rr_func_cmpp_eq_inst24_0_stage_10_o0 & phasebus_0;
  assign and2n_inst269_o0 = rr_func_cmpp_eq_inst23_stage_10_o0 & phasebus_0;
  assign and2n_inst270_o0 = rr_func_cmpp_eq_inst19_stage_10_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst19(
                      .enable0(or2n_inst59_o0),
                      .enable1(and2n_inst272_o0),
                      .i0(select_2_1_wn_inst20_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst19_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst20(
                      .enable0(and2n_inst267_o0),
                      .enable1(and2n_inst270_o0),
                      .i0(sext_inst76_o0[1 : 0]),
                      .i1(sext_inst39_o0[1 : 0]),
                      .o0(select_2_1_wn_inst20_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst76(
                      .i0(1'b0),
                      .o0(sext_inst76_o0[1 : 0]));

  assign or3n_inst45_o0 = and2n_inst268_o0 | and2n_inst269_o0 | and2n_inst266_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:69:7  
  sregn_noinitreset #(.width(2))  rr_var_cbarsactive_stage_11(
                      .clk(clk),
                      .enable(and2n_inst274_o0),
                      .i0(select_2_1_wn_inst19_o0[1 : 0]),
                      .o0(rr_var_cbarsactive_stage_11_o0[1 : 0]));

  assign and2n_inst271_o0 = or3n_inst44_o0 & and3n_inst0_o0;
  assign inverter1n_inst33_o0 = ~or2n_inst59_o0;
  assign and2n_inst272_o0 = sig_start & inverter1n_inst33_o0;
  assign or3n_inst46_o0 = and2n_inst266_o0 | and2n_inst267_o0 | and2n_inst268_o0;
  assign or2n_inst63_o0 = and2n_inst269_o0 | and2n_inst270_o0;
  assign or2n_inst64_o0 = or3n_inst46_o0 | or2n_inst63_o0;
  assign inverter1n_inst34_o0 = ~and2n_inst273_o0;
  assign and2n_inst273_o0 = or3n_inst45_o0 & or2n_inst64_o0;
  assign and2n_inst274_o0 = and2n_inst271_o0 & inverter1n_inst34_o0;
  assign or2n_inst65_o0 = and2n_inst275_o0 | and2n_inst276_o0;
  assign or3n_inst47_o0 = and2n_inst276_o0 | sig_start | phasebus_0;
  assign inverter1n_inst35_o0 = ~and2n_inst276_o0;
  assign and2n_inst275_o0 = inverter1n_inst35_o0 & phasebus_0;
  assign and2n_inst276_o0 = rr_func_cmpp_eq_inst23_0_stage_10_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(2))  select_2_1_wn_inst21(
                      .enable0(or2n_inst65_o0),
                      .enable1(and2n_inst278_o0),
                      .i0(datamerge_select_2_1_wn_inst33_o0[1 : 0]),
                      .i1(2'b00),
                      .o0(select_2_1_wn_inst21_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:69:24  
  sregn_noinitreset #(.width(2))  rr_var_castactive_stage_11(
                      .clk(clk),
                      .enable(and2n_inst280_o0),
                      .i0(select_2_1_wn_inst21_o0[1 : 0]),
                      .o0(rr_var_castactive_stage_11_o0[1 : 0]));

  assign and2n_inst277_o0 = or3n_inst47_o0 & and3n_inst0_o0;
  assign inverter1n_inst36_o0 = ~or2n_inst65_o0;
  assign and2n_inst278_o0 = sig_start & inverter1n_inst36_o0;
  assign or2n_inst67_o0 = and2n_inst275_o0 | and2n_inst276_o0;
  assign nor2n_inst2_o0 = ~(and3n_inst3_o0 | and2n_inst279_o0);
  assign and3n_inst3_o0 = nor2n_inst7_o0 & and2n_inst276_o0 & or2n_inst67_o0;
  assign and2n_inst279_o0 = and2n_inst275_o0 & or2n_inst67_o0;
  assign and2n_inst280_o0 = and2n_inst277_o0 & nor2n_inst2_o0;
  assign and2n_inst281_o0 = cmpp_eq_inst23_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst282_o0),
                      .i0(cmpp_eq_inst23_o0),
                      .o0(rr_func_cmpp_eq_inst23_stage_8_o0));

  assign and2n_inst282_o0 = and2n_inst281_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst283_o0),
                      .i0(rr_func_cmpp_eq_inst23_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst23_stage_9_o0));

  assign and2n_inst283_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst284_o0),
                      .i0(rr_func_cmpp_eq_inst23_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst23_stage_10_o0));

  assign and2n_inst284_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst285_o0),
                      .i0(rr_func_cmpp_eq_inst23_stage_10_o0),
                      .o0(rr_func_cmpp_eq_inst23_stage_11_o0));

  assign and2n_inst285_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst286_o0 = cmpp_eq_inst23_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_0_stage_8(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst287_o0),
                      .i0(cmpp_eq_inst23_o1),
                      .o0(rr_func_cmpp_eq_inst23_0_stage_8_o0));

  assign and2n_inst287_o0 = and2n_inst286_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_0_stage_9(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst288_o0),
                      .i0(rr_func_cmpp_eq_inst23_0_stage_8_o0),
                      .o0(rr_func_cmpp_eq_inst23_0_stage_9_o0));

  assign and2n_inst288_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:115:10  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst23_0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst289_o0),
                      .i0(rr_func_cmpp_eq_inst23_0_stage_9_o0),
                      .o0(rr_func_cmpp_eq_inst23_0_stage_10_o0));

  assign and2n_inst289_o0 = phasebus_0 & and3n_inst0_o0;
  assign or3n_inst48_o0 = and2n_inst290_o0 | and2n_inst291_o0 | and2n_inst292_o0;
  assign or2n_inst68_o0 = or3n_inst48_o0 | and2n_inst293_o0;
  assign or3n_inst49_o0 = and2n_inst293_o0 | and2n_inst291_o0 | and2n_inst292_o0;
  assign or3n_inst50_o0 = or3n_inst49_o0 | sig_start | phasebus_0;
  assign inverter1n_inst37_o0 = ~or3n_inst49_o0;
  assign and2n_inst290_o0 = inverter1n_inst37_o0 & phasebus_0;
  assign and2n_inst291_o0 = rr_func_cmpp_eq_inst20_0_stage_7_o0 & phasebus_0;
  assign and2n_inst292_o0 = rr_func_cmpp_eq_inst21_stage_7_o0 & phasebus_0;
  assign and2n_inst293_o0 = rr_func_cmpp_eq_inst21_0_stage_7_o0 & phasebus_0;

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst22(
                      .enable0(or2n_inst68_o0),
                      .enable1(and2n_inst295_o0),
                      .i0(select_2_1_wn_inst23_o0[11 : 0]),
                      .i1(12'b000000000000),
                      .o0(select_2_1_wn_inst22_o0[11 : 0]));

  select_2_1_wn #(.dwidth(12))  select_2_1_wn_inst23(
                      .enable0(or2n_inst71_o0),
                      .enable1(and2n_inst293_o0),
                      .i0(datamerge_select_2_1_wn_inst32_o0[11 : 0]),
                      .i1(addw_inst2_o0[11 : 0]),
                      .o0(select_2_1_wn_inst23_o0[11 : 0]));

  assign or2n_inst71_o0 = and2n_inst291_o0 | and2n_inst292_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:65:23  
  sregn_noinitreset #(.width(12))  rr_var_ya_1_stage_8(
                      .clk(clk),
                      .enable(and2n_inst297_o0),
                      .i0(select_2_1_wn_inst22_o0[11 : 0]),
                      .o0(rr_var_ya_1_stage_8_o0[11 : 0]));

  assign and2n_inst294_o0 = or3n_inst50_o0 & and3n_inst0_o0;
  assign inverter1n_inst38_o0 = ~or2n_inst68_o0;
  assign and2n_inst295_o0 = sig_start & inverter1n_inst38_o0;
  assign or3n_inst51_o0 = and2n_inst290_o0 | and2n_inst291_o0 | and2n_inst292_o0;
  assign or2n_inst72_o0 = or3n_inst51_o0 | and2n_inst293_o0;
  assign inverter1n_inst39_o0 = ~and2n_inst296_o0;
  assign and2n_inst296_o0 = and2n_inst290_o0 & or2n_inst72_o0;
  assign and2n_inst297_o0 = and2n_inst294_o0 & inverter1n_inst39_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:65:23  
  sregn_noinitreset #(.width(12))  rr_var_ya_1_stage_9(
                      .clk(clk),
                      .enable(and2n_inst298_o0),
                      .i0(rr_var_ya_1_stage_8_o0[11 : 0]),
                      .o0(rr_var_ya_1_stage_9_o0[11 : 0]));

  assign and2n_inst298_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:65:23  
  sregn_noinitreset #(.width(12))  rr_var_ya_1_stage_10(
                      .clk(clk),
                      .enable(and2n_inst299_o0),
                      .i0(rr_var_ya_1_stage_9_o0[11 : 0]),
                      .o0(rr_var_ya_1_stage_10_o0[11 : 0]));

  assign and2n_inst299_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst300_o0 = shrkw_inst2_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:117:31  
  sregn_noinitreset #(.width(30))  rr_func_shrkw_inst2_stage_9(
                      .clk(clk),
                      .enable(and2n_inst301_o0),
                      .i0(shrkw_inst2_o0[29 : 0]),
                      .o0(rr_func_shrkw_inst2_stage_9_o0[29 : 0]));

  assign and2n_inst301_o0 = and2n_inst300_o0 & and3n_inst0_o0;
  assign and2n_inst302_o0 = cmpp_eq_inst24_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:117:17  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst24_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst303_o0),
                      .i0(cmpp_eq_inst24_o0),
                      .o0(rr_func_cmpp_eq_inst24_stage_10_o0));

  assign and2n_inst303_o0 = and2n_inst302_o0 & and3n_inst0_o0;
  assign and2n_inst304_o0 = cmpp_eq_inst24_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:117:17  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst24_0_stage_10(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst305_o0),
                      .i0(cmpp_eq_inst24_o1),
                      .o0(rr_func_cmpp_eq_inst24_0_stage_10_o0));

  assign and2n_inst305_o0 = and2n_inst304_o0 & and3n_inst0_o0;
  assign and2n_inst306_o0 = cmpp_neq_inst1_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:122:6  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst1_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst307_o0),
                      .i0(cmpp_neq_inst1_o0),
                      .o0(rr_func_cmpp_neq_inst1_stage_11_o0));

  assign and2n_inst307_o0 = and2n_inst306_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:122:6  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst1_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst308_o0),
                      .i0(rr_func_cmpp_neq_inst1_stage_11_o0),
                      .o0(rr_func_cmpp_neq_inst1_stage_12_o0));

  assign and2n_inst308_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst309_o0 = cmpp_neq_inst1_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:122:6  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst1_0_stage_11(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst310_o0),
                      .i0(cmpp_neq_inst1_o1),
                      .o0(rr_func_cmpp_neq_inst1_0_stage_11_o0));

  assign and2n_inst310_o0 = and2n_inst309_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:122:6  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst1_0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst311_o0),
                      .i0(rr_func_cmpp_neq_inst1_0_stage_11_o0),
                      .o0(rr_func_cmpp_neq_inst1_0_stage_12_o0));

  assign and2n_inst311_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst312_o0 = cmpp_neq_inst2_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:123:7  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst2_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst313_o0),
                      .i0(cmpp_neq_inst2_o0),
                      .o0(rr_func_cmpp_neq_inst2_stage_12_o0));

  assign and2n_inst313_o0 = and2n_inst312_o0 & and3n_inst0_o0;
  assign and2n_inst314_o0 = cmpp_neq_inst2_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:123:7  
  sregn_noinit #(.width(1))  rr_func_cmpp_neq_inst2_0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst315_o0),
                      .i0(cmpp_neq_inst2_o1),
                      .o0(rr_func_cmpp_neq_inst2_0_stage_12_o0));

  assign and2n_inst315_o0 = and2n_inst314_o0 & and3n_inst0_o0;
  assign and2n_inst316_o0 = cmpp_eq_inst8_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:19  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst8_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst317_o0),
                      .i0(cmpp_eq_inst8_o0),
                      .o0(rr_func_cmpp_eq_inst8_stage_12_o0));

  assign and2n_inst317_o0 = and2n_inst316_o0 & and3n_inst0_o0;
  assign and2n_inst318_o0 = cmpp_eq_inst8_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:19  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst8_0_stage_12(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst319_o0),
                      .i0(cmpp_eq_inst8_o1),
                      .o0(rr_func_cmpp_eq_inst8_0_stage_12_o0));

  assign and2n_inst319_o0 = and2n_inst318_o0 & and3n_inst0_o0;
  assign and2n_inst320_o0 = cmpr_neq_inst5_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:124:31  
  sregn_noinitreset #(.width(2))  rr_func_cmpr_neq_inst5_stage_12(
                      .clk(clk),
                      .enable(and2n_inst321_o0),
                      .i0(cmpr_neq_inst5_o0[1 : 0]),
                      .o0(rr_func_cmpr_neq_inst5_stage_12_o0[1 : 0]));

  assign and2n_inst321_o0 = and2n_inst320_o0 & and3n_inst0_o0;
  assign and2n_inst322_o0 = cmpr_neq_inst6_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:125:31  
  sregn_noinitreset #(.width(2))  rr_func_cmpr_neq_inst6_stage_12(
                      .clk(clk),
                      .enable(and2n_inst323_o0),
                      .i0(cmpr_neq_inst6_o0[1 : 0]),
                      .o0(rr_func_cmpr_neq_inst6_stage_12_o0[1 : 0]));

  assign and2n_inst323_o0 = and2n_inst322_o0 & and3n_inst0_o0;
  assign and2n_inst324_o0 = addw_inst10_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:18  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst10_stage_0(
                      .clk(clk),
                      .enable(and2n_inst325_o0),
                      .i0(addw_inst10_o0[31 : 0]),
                      .o0(rr_func_addw_inst10_stage_0_o0[31 : 0]));

  assign and2n_inst325_o0 = and2n_inst324_o0 & and3n_inst0_o0;
  assign and2n_inst326_o0 = addw_inst11_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:38  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst11_stage_1(
                      .clk(clk),
                      .enable(and2n_inst327_o0),
                      .i0(addw_inst11_o0[31 : 0]),
                      .o0(rr_func_addw_inst11_stage_1_o0[31 : 0]));

  assign and2n_inst327_o0 = and2n_inst326_o0 & and3n_inst0_o0;
  assign and2n_inst328_o0 = addsubw_inst0_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:48  
  sregn_noinitreset #(.width(32))  rr_func_addsubw_inst0_stage_2(
                      .clk(clk),
                      .enable(and2n_inst329_o0),
                      .i0(addsubw_inst0_o0[31 : 0]),
                      .o0(rr_func_addsubw_inst0_stage_2_o0[31 : 0]));

  assign and2n_inst329_o0 = and2n_inst328_o0 & and3n_inst0_o0;
  assign and2n_inst330_o0 = cmpp_eq_inst20_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst331_o0),
                      .i0(cmpp_eq_inst20_o0),
                      .o0(rr_func_cmpp_eq_inst20_stage_3_o0));

  assign and2n_inst331_o0 = and2n_inst330_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst332_o0),
                      .i0(rr_func_cmpp_eq_inst20_stage_3_o0),
                      .o0(rr_func_cmpp_eq_inst20_stage_4_o0));

  assign and2n_inst332_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst333_o0),
                      .i0(rr_func_cmpp_eq_inst20_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst20_stage_5_o0));

  assign and2n_inst333_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst334_o0),
                      .i0(rr_func_cmpp_eq_inst20_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst20_stage_6_o0));

  assign and2n_inst334_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst335_o0 = cmpp_eq_inst20_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_0_stage_3(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst336_o0),
                      .i0(cmpp_eq_inst20_o1),
                      .o0(rr_func_cmpp_eq_inst20_0_stage_3_o0));

  assign and2n_inst336_o0 = and2n_inst335_o0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_0_stage_4(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst337_o0),
                      .i0(rr_func_cmpp_eq_inst20_0_stage_3_o0),
                      .o0(rr_func_cmpp_eq_inst20_0_stage_4_o0));

  assign and2n_inst337_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_0_stage_5(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst338_o0),
                      .i0(rr_func_cmpp_eq_inst20_0_stage_4_o0),
                      .o0(rr_func_cmpp_eq_inst20_0_stage_5_o0));

  assign and2n_inst338_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_0_stage_6(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst339_o0),
                      .i0(rr_func_cmpp_eq_inst20_0_stage_5_o0),
                      .o0(rr_func_cmpp_eq_inst20_0_stage_6_o0));

  assign and2n_inst339_o0 = phasebus_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:141:8  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst20_0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst340_o0),
                      .i0(rr_func_cmpp_eq_inst20_0_stage_6_o0),
                      .o0(rr_func_cmpp_eq_inst20_0_stage_7_o0));

  assign and2n_inst340_o0 = phasebus_0 & and3n_inst0_o0;
  assign and2n_inst341_o0 = addw_inst12_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:19  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst12_stage_4(
                      .clk(clk),
                      .enable(and2n_inst342_o0),
                      .i0(addw_inst12_o0[31 : 0]),
                      .o0(rr_func_addw_inst12_stage_4_o0[31 : 0]));

  assign and2n_inst342_o0 = and2n_inst341_o0 & and3n_inst0_o0;
  assign and2n_inst343_o0 = addw_inst13_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:39  
  sregn_noinitreset #(.width(32))  rr_func_addw_inst13_stage_5(
                      .clk(clk),
                      .enable(and2n_inst344_o0),
                      .i0(addw_inst13_o0[31 : 0]),
                      .o0(rr_func_addw_inst13_stage_5_o0[31 : 0]));

  assign and2n_inst344_o0 = and2n_inst343_o0 & and3n_inst0_o0;
  assign and2n_inst345_o0 = addsubw_inst1_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:49  
  sregn_noinitreset #(.width(32))  rr_func_addsubw_inst1_stage_6(
                      .clk(clk),
                      .enable(and2n_inst346_o0),
                      .i0(addsubw_inst1_o0[31 : 0]),
                      .o0(rr_func_addsubw_inst1_stage_6_o0[31 : 0]));

  assign and2n_inst346_o0 = and2n_inst345_o0 & and3n_inst0_o0;
  assign and2n_inst347_o0 = cmpp_eq_inst21_o0_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:9  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst21_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst348_o0),
                      .i0(cmpp_eq_inst21_o0),
                      .o0(rr_func_cmpp_eq_inst21_stage_7_o0));

  assign and2n_inst348_o0 = and2n_inst347_o0 & and3n_inst0_o0;
  assign and2n_inst349_o0 = cmpp_eq_inst21_o1_enable & phasebus_0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:142:9  
  sregn_noinit #(.width(1))  rr_func_cmpp_eq_inst21_0_stage_7(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst350_o0),
                      .i0(cmpp_eq_inst21_o1),
                      .o0(rr_func_cmpp_eq_inst21_0_stage_7_o0));

  assign and2n_inst350_o0 = and2n_inst349_o0 & and3n_inst0_o0;

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst24(
                      .enable0(cmpp_eq_inst2_o0),
                      .enable1(cmpp_eq_inst2_o1),
                      .i0(sext_inst77_o0[1 : 0]),
                      .i1(sext_inst17_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst24_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst77(
                      .i0(1'b0),
                      .o0(sext_inst77_o0[1 : 0]));

  select_2_1_wn #(.dwidth(1))  datamerge_select_2_1_wn_inst25(
                      .enable0(rr_func_cmpp_eq_inst0_stage_6_o0),
                      .enable1(rr_func_cmpp_eq_inst12_stage_6_o0),
                      .i0(datamerge_select_2_1_wn_inst24_o0[0]),
                      .i1(datamerge_select_2_1_wn_inst26_o0[0]),
                      .o0(datamerge_select_2_1_wn_inst25_o0));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst26(
                      .enable0(cmpp_eq_inst3_o0),
                      .enable1(cmpp_eq_inst3_o1),
                      .i0(sext_inst18_o0[1 : 0]),
                      .i1(sext_inst78_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst26_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst78(
                      .i0(1'b0),
                      .o0(sext_inst78_o0[1 : 0]));

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst2(
                      .enable0(rr_func_cmpp_eq_inst13_stage_12_o0),
                      .enable1(or3n_inst53_o0),
                      .enable2(rr_func_cmpp_eq_inst14_stage_12_o0),
                      .i0(sext_inst19_o0[1 : 0]),
                      .i1(rr_var_hactive_stage_13_o0[1 : 0]),
                      .i2(sext_inst79_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst2_o0[1 : 0]));

  assign or3n_inst53_o0 = rr_func_cmpp_eq_inst12_stage_12_o0 | rr_func_cmpp_eq_inst0_stage_12_o0 | rr_func_cmpp_eq_inst14_0_stage_12_o0;

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst79(
                      .i0(1'b0),
                      .o0(sext_inst79_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst27(
                      .enable0(cmpp_eq_inst4_o0),
                      .enable1(cmpp_eq_inst4_o1),
                      .i0(sext_inst80_o0[1 : 0]),
                      .i1(sext_inst21_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst27_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst80(
                      .i0(1'b0),
                      .o0(sext_inst80_o0[1 : 0]));

  select_3_1_wn #(.dwidth(1))  datamerge_select_3_1_wn_inst3(
                      .enable0(rr_func_cmpp_eq_inst1_stage_12_o0),
                      .enable1(rr_func_cmpp_eq_inst15_stage_12_o0),
                      .enable2(nor2n_inst4_o0),
                      .i0(datamerge_select_2_1_wn_inst27_o0[0]),
                      .i1(datamerge_select_2_1_wn_inst29_o0[0]),
                      .i2(rr_var_dvi_ds_s_vs_stage_12_o0),
                      .o0(datamerge_select_3_1_wn_inst3_o0));

  select_2_1_wn #(.dwidth(1))  datamerge_select_2_1_wn_inst28(
                      .enable0(rr_func_cmpp_eq_inst1_stage_12_o0),
                      .enable1(rr_func_cmpp_eq_inst15_stage_12_o0),
                      .i0(datamerge_select_2_1_wn_inst27_o0[0]),
                      .i1(datamerge_select_2_1_wn_inst29_o0[0]),
                      .o0(datamerge_select_2_1_wn_inst28_o0));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst29(
                      .enable0(cmpp_eq_inst5_o0),
                      .enable1(cmpp_eq_inst5_o1),
                      .i0(sext_inst22_o0[1 : 0]),
                      .i1(sext_inst81_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst29_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst81(
                      .i0(1'b0),
                      .o0(sext_inst81_o0[1 : 0]));

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst4(
                      .enable0(rr_func_cmpp_eq_inst16_stage_12_o0),
                      .enable1(or3n_inst56_o0),
                      .enable2(rr_func_cmpp_eq_inst17_stage_12_o0),
                      .i0(sext_inst23_o0[1 : 0]),
                      .i1(rr_var_vactive_stage_13_o0[1 : 0]),
                      .i2(sext_inst82_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst4_o0[1 : 0]));

  assign or3n_inst56_o0 = rr_func_cmpp_eq_inst15_stage_12_o0 | rr_func_cmpp_eq_inst1_stage_12_o0 | rr_func_cmpp_eq_inst17_0_stage_12_o0;

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst82(
                      .i0(1'b0),
                      .o0(sext_inst82_o0[1 : 0]));

  select_2_1_wn #(.dwidth(12))  datamerge_select_2_1_wn_inst30(
                      .enable0(rr_func_cmpp_eq_inst18_stage_4_o0),
                      .enable1(inverter1n_inst40_o0),
                      .i0(sext_inst83_o0[11 : 0]),
                      .i1(rr_var_xa_stage_4_o0[11 : 0]),
                      .o0(datamerge_select_2_1_wn_inst30_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst83(
                      .i0(1'b0),
                      .o0(sext_inst83_o0[11 : 0]));

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst5(
                      .enable0(rr_func_cmpp_eq_inst18_stage_11_o0),
                      .enable1(rr_func_cmpp_eq_inst22_0_stage_11_o0),
                      .enable2(rr_func_cmpp_eq_inst22_stage_11_o0),
                      .i0(sext_inst24_o0[1 : 0]),
                      .i1(rr_var_bactive_stage_12_o0[1 : 0]),
                      .i2(rr_func_moveii_inst40_stage_11_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst5_o0[1 : 0]));

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst6(
                      .enable0(rr_func_cmpp_eq_inst18_stage_11_o0),
                      .enable1(or2n_inst80_o0),
                      .enable2(cmpp_eq_inst6_o0),
                      .i0(sext_inst25_o0[1 : 0]),
                      .i1(rr_var_gactive_stage_12_o0[1 : 0]),
                      .i2(cmpr_eq_inst2_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst6_o0[1 : 0]));

  assign or2n_inst80_o0 = cmpp_eq_inst6_o1 | rr_func_cmpp_eq_inst22_0_stage_11_o0;

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst7(
                      .enable0(rr_func_cmpp_eq_inst18_stage_11_o0),
                      .enable1(or2n_inst81_o0),
                      .enable2(cmpp_eq_inst7_o0),
                      .i0(sext_inst26_o0[1 : 0]),
                      .i1(rr_var_ractive_stage_12_o0[1 : 0]),
                      .i2(cmpr_eq_inst3_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst7_o0[1 : 0]));

  assign or2n_inst81_o0 = cmpp_eq_inst7_o1 | rr_func_cmpp_eq_inst22_0_stage_11_o0;

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst31(
                      .enable0(rr_func_cmpp_neq_inst0_stage_11_o0),
                      .enable1(cmpr_eq_inst1_o0_enable),
                      .i0(rr_func_moveii_inst40_stage_11_o0[1 : 0]),
                      .i1(cmpr_eq_inst1_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst31_o0[1 : 0]));

  select_2_1_wn #(.dwidth(12))  datamerge_select_2_1_wn_inst32(
                      .enable0(rr_func_cmpp_eq_inst19_stage_7_o0),
                      .enable1(rr_func_cmpp_eq_inst19_0_stage_7_o0),
                      .i0(sext_inst84_o0[11 : 0]),
                      .i1(rr_var_ya_1_stage_8_o0[11 : 0]),
                      .o0(datamerge_select_2_1_wn_inst32_o0[11 : 0]));

  sext #(.inwidth(1), .outwidth(12), .signedflag(0))  sext_inst84(
                      .i0(1'b0),
                      .o0(sext_inst84_o0[11 : 0]));

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst8(
                      .enable0(rr_func_cmpp_eq_inst19_stage_10_o0),
                      .enable1(or2n_inst84_o0),
                      .enable2(rr_func_cmpp_eq_inst24_stage_10_o0),
                      .i0(sext_inst39_o0[1 : 0]),
                      .i1(rr_var_cbarsactive_stage_11_o0[1 : 0]),
                      .i2(sext_inst85_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst8_o0[1 : 0]));

  assign or2n_inst84_o0 = rr_func_cmpp_eq_inst23_stage_10_o0 | rr_func_cmpp_eq_inst24_0_stage_10_o0;

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst85(
                      .i0(1'b0),
                      .o0(sext_inst85_o0[1 : 0]));

  select_3_1_wn #(.dwidth(2))  datamerge_select_3_1_wn_inst9(
                      .enable0(rr_func_cmpp_eq_inst19_stage_11_o0),
                      .enable1(rr_func_cmpp_eq_inst23_stage_11_o0),
                      .enable2(nor2n_inst6_o0),
                      .i0(sext_inst86_o0[1 : 0]),
                      .i1(sext_inst40_o0[1 : 0]),
                      .i2(rr_var_castactive_stage_11_o0[1 : 0]),
                      .o0(datamerge_select_3_1_wn_inst9_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst86(
                      .i0(1'b0),
                      .o0(sext_inst86_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst33(
                      .enable0(rr_func_cmpp_eq_inst19_stage_11_o0),
                      .enable1(rr_func_cmpp_eq_inst23_stage_11_o0),
                      .i0(sext_inst87_o0[1 : 0]),
                      .i1(sext_inst40_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst33_o0[1 : 0]));

  sext #(.inwidth(1), .outwidth(2), .signedflag(1))  sext_inst87(
                      .i0(1'b0),
                      .o0(sext_inst87_o0[1 : 0]));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst34(
                      .enable0(rr_func_cmpp_eq_inst8_stage_12_o0),
                      .enable1(cmpr_eq_inst4_o0_enable),
                      .i0(cmpr_neq_inst4_o0[1 : 0]),
                      .i1(cmpr_eq_inst4_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst34_o0[1 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst35(
                      .enable0(cmpp_eq_inst9_o0),
                      .enable1(cmpp_eq_inst9_o1),
                      .i0(sext_inst48_o0[8 : 0]),
                      .i1(sext_inst88_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst35_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst88(
                      .i0(1'b0),
                      .o0(sext_inst88_o0[8 : 0]));

  select_3_1_wn #(.dwidth(8))  datamerge_select_3_1_wn_inst10(
                      .enable0(rr_func_cmpp_neq_inst2_stage_12_o0),
                      .enable1(rr_func_cmpp_neq_inst2_0_stage_12_o0),
                      .enable2(rr_func_cmpp_neq_inst1_0_stage_12_o0),
                      .i0(datamerge_select_2_1_wn_inst35_o0[7 : 0]),
                      .i1(datamerge_select_2_1_wn_inst38_o0[7 : 0]),
                      .i2(datamerge_select_2_1_wn_inst42_o0[7 : 0]),
                      .o0(datamerge_select_3_1_wn_inst10_o0[7 : 0]));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst36(
                      .enable0(rr_func_cmpp_eq_inst8_stage_12_o0),
                      .enable1(cmpr_eq_inst5_o0_enable),
                      .i0(cmpr_neq_inst4_o0[1 : 0]),
                      .i1(cmpr_eq_inst5_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst36_o0[1 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst37(
                      .enable0(cmpp_eq_inst10_o0),
                      .enable1(cmpp_eq_inst10_o1),
                      .i0(sext_inst52_o0[8 : 0]),
                      .i1(sext_inst89_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst37_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst89(
                      .i0(1'b0),
                      .o0(sext_inst89_o0[8 : 0]));

  select_3_1_wn #(.dwidth(8))  datamerge_select_3_1_wn_inst11(
                      .enable0(rr_func_cmpp_neq_inst2_stage_12_o0),
                      .enable1(rr_func_cmpp_neq_inst2_0_stage_12_o0),
                      .enable2(rr_func_cmpp_neq_inst1_0_stage_12_o0),
                      .i0(datamerge_select_2_1_wn_inst37_o0[7 : 0]),
                      .i1(datamerge_select_2_1_wn_inst39_o0[7 : 0]),
                      .i2(datamerge_select_2_1_wn_inst43_o0[7 : 0]),
                      .o0(datamerge_select_3_1_wn_inst11_o0[7 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst38(
                      .enable0(cmpp_neq_inst3_o0),
                      .enable1(cmpp_neq_inst3_o1),
                      .i0(sext_inst54_o0[8 : 0]),
                      .i1(sext_inst90_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst38_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst90(
                      .i0(1'b0),
                      .o0(sext_inst90_o0[8 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst39(
                      .enable0(cmpp_neq_inst4_o0),
                      .enable1(cmpp_neq_inst4_o1),
                      .i0(sext_inst56_o0[8 : 0]),
                      .i1(sext_inst91_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst39_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst91(
                      .i0(1'b0),
                      .o0(sext_inst91_o0[8 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst40(
                      .enable0(cmpp_neq_inst5_o0),
                      .enable1(cmpp_neq_inst5_o1),
                      .i0(sext_inst58_o0[8 : 0]),
                      .i1(sext_inst92_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst40_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst92(
                      .i0(1'b0),
                      .o0(sext_inst92_o0[8 : 0]));

  select_2_1_wn #(.dwidth(8))  datamerge_select_2_1_wn_inst41(
                      .enable0(rr_func_cmpp_neq_inst1_stage_12_o0),
                      .enable1(rr_func_cmpp_neq_inst1_0_stage_12_o0),
                      .i0(datamerge_select_2_1_wn_inst40_o0[7 : 0]),
                      .i1(datamerge_select_2_1_wn_inst44_o0[7 : 0]),
                      .o0(datamerge_select_2_1_wn_inst41_o0[7 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst42(
                      .enable0(cmpp_neq_inst6_o0),
                      .enable1(cmpp_neq_inst6_o1),
                      .i0(sext_inst60_o0[8 : 0]),
                      .i1(sext_inst93_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst42_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst93(
                      .i0(1'b0),
                      .o0(sext_inst93_o0[8 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst43(
                      .enable0(cmpp_neq_inst6_o0),
                      .enable1(cmpp_neq_inst6_o1),
                      .i0(sext_inst61_o0[8 : 0]),
                      .i1(sext_inst94_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst43_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst94(
                      .i0(1'b0),
                      .o0(sext_inst94_o0[8 : 0]));

  select_2_1_wn #(.dwidth(9))  datamerge_select_2_1_wn_inst44(
                      .enable0(cmpp_neq_inst6_o0),
                      .enable1(cmpp_neq_inst6_o1),
                      .i0(sext_inst62_o0[8 : 0]),
                      .i1(sext_inst95_o0[8 : 0]),
                      .o0(datamerge_select_2_1_wn_inst44_o0[8 : 0]));

  sext #(.inwidth(1), .outwidth(9), .signedflag(1))  sext_inst95(
                      .i0(1'b0),
                      .o0(sext_inst95_o0[8 : 0]));

  select_2_1_wn #(.dwidth(2))  datamerge_select_2_1_wn_inst45(
                      .enable0(cmpp_eq_inst11_o0),
                      .enable1(cmpr_neq_inst8_o0_enable),
                      .i0(cmpr_neq_inst7_o0[1 : 0]),
                      .i1(cmpr_neq_inst8_o0[1 : 0]),
                      .o0(datamerge_select_2_1_wn_inst45_o0[1 : 0]));

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:56:14  
  sregn_noinit #(.width(1))  sr_var_hsync(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst351_o0),
                      .i0(sig_lid_rawdatain_hsync_0_0),
                      .o0(sr_var_hsync_o0));

  assign and2n_inst351_o0 = sig_lien_rawdatain_hsync_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:54:14  
  sregn_noinitreset #(.width(32))  sr_var_hblank(
                      .clk(clk),
                      .enable(and2n_inst352_o0),
                      .i0(sig_lid_rawdatain_hblank_0_0[31 : 0]),
                      .o0(sr_var_hblank_o0[31 : 0]));

  assign and2n_inst352_o0 = sig_lien_rawdatain_hblank_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:55:14  
  sregn_noinitreset #(.width(32))  sr_var_hbporch(
                      .clk(clk),
                      .enable(and2n_inst353_o0),
                      .i0(sig_lid_rawdatain_hbporch_0_0[31 : 0]),
                      .o0(sr_var_hbporch_o0[31 : 0]));

  assign and2n_inst353_o0 = sig_lien_rawdatain_hbporch_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:52:14  
  sregn_noinitreset #(.width(32))  sr_var_hactive_1(
                      .clk(clk),
                      .enable(and2n_inst354_o0),
                      .i0(sig_lid_rawdatain_hactive_0_0[31 : 0]),
                      .o0(sr_var_hactive_1_o0[31 : 0]));

  assign and2n_inst354_o0 = sig_lien_rawdatain_hactive_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:57:14  
  sregn_noinit #(.width(1))  sr_var_vsync(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst355_o0),
                      .i0(sig_lid_rawdatain_vsync_0_0),
                      .o0(sr_var_vsync_o0));

  assign and2n_inst355_o0 = sig_lien_rawdatain_vsync_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:50:14  
  sregn_noinitreset #(.width(32))  sr_var_vblank(
                      .clk(clk),
                      .enable(and2n_inst356_o0),
                      .i0(sig_lid_rawdatain_vblank_0_0[31 : 0]),
                      .o0(sr_var_vblank_o0[31 : 0]));

  assign and2n_inst356_o0 = sig_lien_rawdatain_vblank_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:51:14  
  sregn_noinitreset #(.width(32))  sr_var_vbporch(
                      .clk(clk),
                      .enable(and2n_inst357_o0),
                      .i0(sig_lid_rawdatain_vbporch_0_0[31 : 0]),
                      .o0(sr_var_vbporch_o0[31 : 0]));

  assign and2n_inst357_o0 = sig_lien_rawdatain_vbporch_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:48:14  
  sregn_noinitreset #(.width(32))  sr_var_vactive_1(
                      .clk(clk),
                      .enable(and2n_inst358_o0),
                      .i0(sig_lid_rawdatain_vactive_0_0[31 : 0]),
                      .o0(sr_var_vactive_1_o0[31 : 0]));

  assign and2n_inst358_o0 = sig_lien_rawdatain_vactive_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:53:14  
  sregn_noinitreset #(.width(32))  sr_var_hfporch(
                      .clk(clk),
                      .enable(and2n_inst359_o0),
                      .i0(sig_lid_rawdatain_hfporch_0_0[31 : 0]),
                      .o0(sr_var_hfporch_o0[31 : 0]));

  assign and2n_inst359_o0 = sig_lien_rawdatain_hfporch_0_0 & and3n_inst0_o0;

  // dvi_interface/test_pattern_generator/test_pattern_generator.cpp:49:14  
  sregn_noinitreset #(.width(32))  sr_var_vfporch(
                      .clk(clk),
                      .enable(and2n_inst360_o0),
                      .i0(sig_lid_rawdatain_vfporch_0_0[31 : 0]),
                      .o0(sr_var_vfporch_o0[31 : 0]));

  assign and2n_inst360_o0 = sig_lien_rawdatain_vfporch_0_0 & and3n_inst0_o0;

  sregn_noinit #(.width(1))  sr_var_loopcounter(
                      .clk(clk),
                      .reset(reset),
                      .enable(and2n_inst361_o0),
                      .i0(1'b1),
                      .o0(sr_var_loopcounter_o0));

  assign and2n_inst361_o0 = sig_start & and3n_inst0_o0;
  assign nor2n_inst3_o0 = ~(rr_func_cmpp_eq_inst0_stage_6_o0 | rr_func_cmpp_eq_inst12_stage_6_o0);
  assign nor2n_inst4_o0 = ~(rr_func_cmpp_eq_inst1_stage_12_o0 | rr_func_cmpp_eq_inst15_stage_12_o0);
  assign nor2n_inst5_o0 = ~(rr_func_cmpp_eq_inst1_stage_12_o0 | rr_func_cmpp_eq_inst15_stage_12_o0);
  assign inverter1n_inst40_o0 = ~rr_func_cmpp_eq_inst18_stage_4_o0;
  assign nor3n_inst0_o0 = ~(rr_func_cmpp_eq_inst18_stage_11_o0 | rr_func_cmpp_eq_inst22_0_stage_11_o0 | rr_func_cmpp_eq_inst22_stage_11_o0);
  assign nor2n_inst6_o0 = ~(rr_func_cmpp_eq_inst19_stage_11_o0 | rr_func_cmpp_eq_inst23_stage_11_o0);
  assign nor2n_inst7_o0 = ~(rr_func_cmpp_eq_inst19_stage_11_o0 | rr_func_cmpp_eq_inst23_stage_11_o0);
  assign inverter1n_inst41_o0 = ~outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0_stallbar;
  assign inverter1n_inst42_o0 = ~retimed_reg_o0;

  sregn_noinit #(.width(1))  retimed_reg(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .i0(inverter1n_inst41_o0),
                      .o0(retimed_reg_o0));



`ifdef PICO_DUMP_STALL_BREAKUP
// synopsys translate_off
   reg doStallCounting;
   integer stallfptr;
   integer verifyfptr;
   integer count0;
   integer count1;
   integer count2;
   initial begin
           doStallCounting = 0;
           count0 = 1;
           count1 = 1;
           count2 = 1;
    verifyfptr = $fopen("verify.out");
    stallfptr  = $fopen("stalls.out"); end
   always @(posedge enable) begin// Start counting from chip-enable high 
           doStallCounting = 1; // never reset
   end
   always @(posedge clk) begin
      #1;
      if(~outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0.stallbar & doStallCounting) begin
         $fdisplay(verifyfptr,"%d:%m.outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0.stallbar",count0);
	 count0 <= count0 + 1;
         $fdisplay(stallfptr,"%d:%m.outstream_dvi_out_dismantle_test_pattern_generator_wide_ststream0_0_noreset_inst0.stallbar", $stime); end
    end

   always @(posedge clk) begin
      #1;
      if(~stallbar_in & doStallCounting) begin
         $fdisplay(verifyfptr,"%d:%m.stallbar_in",count1);
	 count1 <= count1 + 1;
         $fdisplay(stallfptr,"%d:%m.stallbar_in", $stime); end
    end

   always @(posedge clk) begin
      #1;
      if(~enable & doStallCounting) begin
         $fdisplay(verifyfptr,"%d:%m.enable",count2);
	 count2 <= count2 + 1;
         $fdisplay(stallfptr,"%d:%m.enable", $stime); end
    end

// synopsys translate_on
`endif

endmodule


// vim: tags=./tags_test_pattern_generator_pe_0_v
