/************************************************************************
 *                                                                      *
 * Copyright (c) 2009 Synfora, Inc.  All rights reserved.               *
 *                                                                      *
 * This file contains Confidential Information of Synfora, Inc.         *
 * In addition, certain inventions disclosed in this file may be        *
 * claimed within patents owned or patent applications filed by         *
 * Synfora or third parties.  Any use of Synfora's copyrighted works,   *
 * confidential information, patented inventions, or patent-pending     *
 * inventions is subject to the terms and conditions of your written    *
 * license agreement with Synfora, Inc.                                 *
 * All other use and disclosure is strictly prohibited.                 *
 *                                                                      *
 ************************************************************************/

/* Generated by PICO Extreme FPGA version 09.04 */
/* Target library : xilinx-spartan6-s2 */
/* Target frequency : 100 MHz */

`timescale 1ns / 10 ps

// The following defines named constants used in this file.
`ifdef TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH
`else
`define TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH 0
`endif
// End of definitions of named constants

module test_pattern_generator_ppa(
        clk,
        reset,
        start_task_init,
        start_task_final,
        clear_init_done,
        clear_task_done,
        psw_livein_frames_in_use,
        psw_liveout_frames_in_use,
        psw_released,
        psw_sa_0_stalling,
        psw_busy,
        psw_idle,
        psw_init_done,
        psw_task_done,
        rawdatain_hsync_0,
        rawdatain_hblank_0,
        rawdatain_hbporch_0,
        rawdatain_hactive_0,
        rawdatain_vsync_0,
        rawdatain_vblank_0,
        rawdatain_vbporch_0,
        rawdatain_vactive_0,
        rawdatain_hfporch_0,
        rawdatain_vfporch_0,
        outstream_dvi_out_do_0,
        outstream_dvi_out_req_0,
        outstream_dvi_out_ready_0);

  // Module parameters


  // synopsys template

  // Ports

  input  clk;
  input  reset;
  input  start_task_init;
  input  start_task_final;
  input  clear_init_done;
  input  clear_task_done;
  output [3 : 0] psw_livein_frames_in_use;
  output [3 : 0] psw_liveout_frames_in_use;
  output  psw_released;
  output  psw_sa_0_stalling;
  output  psw_busy;
  output  psw_idle;
  output  psw_init_done;
  output  psw_task_done;
  input  rawdatain_hsync_0;
  input [31 : 0] rawdatain_hblank_0;
  input [31 : 0] rawdatain_hbporch_0;
  input [31 : 0] rawdatain_hactive_0;
  input  rawdatain_vsync_0;
  input [31 : 0] rawdatain_vblank_0;
  input [31 : 0] rawdatain_vbporch_0;
  input [31 : 0] rawdatain_vactive_0;
  input [31 : 0] rawdatain_hfporch_0;
  input [31 : 0] rawdatain_vfporch_0;
  output [26 : 0] outstream_dvi_out_do_0;
  output  outstream_dvi_out_req_0;
  input  outstream_dvi_out_ready_0;

  // Wire/Reg for portformals 

  wire  clk;
  wire  reset;
  wire  start_task_init;
  wire  start_task_final;
  wire  clear_init_done;
  wire  clear_task_done;
  wire [3 : 0] psw_livein_frames_in_use;
  wire [3 : 0] psw_liveout_frames_in_use;
  wire  psw_released;
  wire  psw_sa_0_stalling;
  wire  psw_busy;
  wire  psw_idle;
  wire  psw_init_done;
  wire  psw_task_done;
  wire  rawdatain_hsync_0;
  wire [31 : 0] rawdatain_hblank_0;
  wire [31 : 0] rawdatain_hbporch_0;
  wire [31 : 0] rawdatain_hactive_0;
  wire  rawdatain_vsync_0;
  wire [31 : 0] rawdatain_vblank_0;
  wire [31 : 0] rawdatain_vbporch_0;
  wire [31 : 0] rawdatain_vactive_0;
  wire [31 : 0] rawdatain_hfporch_0;
  wire [31 : 0] rawdatain_vfporch_0;
  wire [26 : 0] outstream_dvi_out_do_0;
  wire  outstream_dvi_out_req_0;
  wire  outstream_dvi_out_ready_0;

  wire [26 : 0] boundary_buf_outstream_dvi_out_dismantle_outdata;
  wire  boundary_buf_outstream_dvi_out_dismantle_store_req;
  wire  sig_outstream_dvi_out_ready_0;
  wire  psw_start_task_init_internal;
  wire  paw_0_status;
  wire  paw_0_err;
  wire  paw_0_busy;
  wire  paw_0_stallbar_out;
  wire [26 : 0] paw_0_outstream_dvi_out_do_0;
  wire  paw_0_outstream_dvi_out_req_0;
  wire  boundary_buf_outstream_dvi_out_dismantle_load_req;
  wire  sig_rawdatain_hsync_0;
  wire [31 : 0] sig_rawdatain_hblank_0;
  wire [31 : 0] sig_rawdatain_hbporch_0;
  wire [31 : 0] sig_rawdatain_hactive_0;
  wire  sig_rawdatain_vsync_0;
  wire [31 : 0] sig_rawdatain_vblank_0;
  wire [31 : 0] sig_rawdatain_vbporch_0;
  wire [31 : 0] sig_rawdatain_vactive_0;
  wire [31 : 0] sig_rawdatain_hfporch_0;
  wire [31 : 0] sig_rawdatain_vfporch_0;
  wire  sig_clk;
  wire  sig_clear_init_done;
  wire  sig_clear_task_done;
  wire [3 : 0] sext_inst0_o0;
  wire [3 : 0] sext_inst1_o0;
  wire  psw_released_internal;
  wire  registered_port_sregn_noinit_inst4_o0;
  wire  psw_busy_internal;
  wire  psw_idle_internal;
  wire  psw_init_done_internal;
  wire  psw_task_done_internal;
  wire  psw_sa_0_stalling_internal;
  wire  reset_pulsereg1_o0;
  wire  inverter1n_inst5_o0;
  wire  reset_pulsereg2_o0;
  wire  sregn_noinit_inst5_dly_o0;
  wire  and2n_inst0_o0;
  wire  inverter1n_inst6_o0;
  wire  and2n_inst2_o0;
  wire  task_done_pulse;
  wire  and2n_inst5_o0;
  wire  inverter1n_inst7_o0;
  wire  psw_livein_frames_in_use_internal;
  wire  psw_liveout_frames_in_use_internal;
  wire  equal_inst0_o0;
  wire  equal_inst1_o0;
  wire  multiloop_rsflipflop_noinit_inst3_q;
  wire  multiloop_rsflipflop_noinit_inst2_q;
  wire  inverter1n_inst8_o0;
  wire  pulsereg_sastatus_0_o0;
  wire  and2n_inst4_o0;
  wire  and2n_inst6_o0;
  wire  and2n_inst7_o0;
  wire  inverter1n_inst10_o0;
  wire  inverter1n_inst11_o0;


  // Signal assignments

  assign outstream_dvi_out_do_0 = boundary_buf_outstream_dvi_out_dismantle_outdata;
  assign outstream_dvi_out_req_0 = boundary_buf_outstream_dvi_out_dismantle_store_req;
  assign sig_outstream_dvi_out_ready_0 = outstream_dvi_out_ready_0;
  assign sig_rawdatain_hsync_0 = rawdatain_hsync_0;
  assign sig_rawdatain_hblank_0 = rawdatain_hblank_0;
  assign sig_rawdatain_hbporch_0 = rawdatain_hbporch_0;
  assign sig_rawdatain_hactive_0 = rawdatain_hactive_0;
  assign sig_rawdatain_vsync_0 = rawdatain_vsync_0;
  assign sig_rawdatain_vblank_0 = rawdatain_vblank_0;
  assign sig_rawdatain_vbporch_0 = rawdatain_vbporch_0;
  assign sig_rawdatain_vactive_0 = rawdatain_vactive_0;
  assign sig_rawdatain_hfporch_0 = rawdatain_hfporch_0;
  assign sig_rawdatain_vfporch_0 = rawdatain_vfporch_0;
  assign sig_clk = clk;
  assign sig_clear_init_done = clear_init_done;
  assign sig_clear_task_done = clear_task_done;
  assign psw_livein_frames_in_use = sext_inst0_o0;
  assign psw_liveout_frames_in_use = sext_inst1_o0;
  assign psw_released = psw_released_internal;
  assign psw_sa_0_stalling = registered_port_sregn_noinit_inst4_o0;
  assign psw_busy = psw_busy_internal;
  assign psw_idle = psw_idle_internal;
  assign psw_init_done = psw_init_done_internal;
  assign psw_task_done = psw_task_done_internal;

  // Basic logic assignments


  // Component port and generic maps / Behavioural code.

  test_pattern_generator_paw_0  paw_0(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .start(psw_start_task_init_internal),
                      .abort(1'b0),
                      .status(paw_0_status),
                      .err(paw_0_err),
                      .stallbar_in(1'b1),
                      .stallbar_out(paw_0_stallbar_out),
                      .busy(paw_0_busy),
                      .outstream_dvi_out_do_0(paw_0_outstream_dvi_out_do_0[26 : 0]),
                      .outstream_dvi_out_req_0(paw_0_outstream_dvi_out_req_0),
                      .outstream_dvi_out_ready_0(boundary_buf_outstream_dvi_out_dismantle_load_req),
                      .rawdatain_0_0(sig_rawdatain_hsync_0),
                      .rawdatainenable_0_0(psw_start_task_init_internal),
                      .rawdatain_1_0(sig_rawdatain_hblank_0[31 : 0]),
                      .rawdatainenable_1_0(psw_start_task_init_internal),
                      .rawdatain_2_0(sig_rawdatain_hbporch_0[31 : 0]),
                      .rawdatainenable_2_0(psw_start_task_init_internal),
                      .rawdatain_3_0(sig_rawdatain_hactive_0[31 : 0]),
                      .rawdatainenable_3_0(psw_start_task_init_internal),
                      .rawdatain_4_0(sig_rawdatain_vsync_0),
                      .rawdatainenable_4_0(psw_start_task_init_internal),
                      .rawdatain_5_0(sig_rawdatain_vblank_0[31 : 0]),
                      .rawdatainenable_5_0(psw_start_task_init_internal),
                      .rawdatain_6_0(sig_rawdatain_vbporch_0[31 : 0]),
                      .rawdatainenable_6_0(psw_start_task_init_internal),
                      .rawdatain_7_0(sig_rawdatain_vactive_0[31 : 0]),
                      .rawdatainenable_7_0(psw_start_task_init_internal),
                      .rawdatain_8_0(sig_rawdatain_hfporch_0[31 : 0]),
                      .rawdatainenable_8_0(psw_start_task_init_internal),
                      .rawdatain_9_0(sig_rawdatain_vfporch_0[31 : 0]),
                      .rawdatainenable_9_0(psw_start_task_init_internal));

  sregn_noinit #(.width(1))  registered_port_sregn_noinit_inst4(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .i0(psw_sa_0_stalling_internal),
                      .o0(registered_port_sregn_noinit_inst4_o0));

  sregn_noinit #(.width(1))  reset_pulsereg1(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .i0(1'b1),
                      .o0(reset_pulsereg1_o0));

  assign inverter1n_inst5_o0 = ~reset_pulsereg1_o0;

  sregn_noinit #(.width(1))  reset_pulsereg2(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .i0(inverter1n_inst5_o0),
                      .o0(reset_pulsereg2_o0));

  assign psw_start_task_init_internal = reset_pulsereg2_o0 | sregn_noinit_inst5_dly_o0;

  rsflipflop_noinit  mlinterface_rsflipflop_noinit_inst0(
                      .clk(clk),
                      .reset(reset),
                      .r(and2n_inst0_o0),
                      .s(psw_start_task_init_internal),
                      .q(psw_init_done_internal));

  assign and2n_inst0_o0 = sig_clear_init_done & inverter1n_inst6_o0;
  assign inverter1n_inst6_o0 = ~psw_start_task_init_internal;

  rsflipflop_noinit  mlinterface_rsflipflop_noinit_inst1(
                      .clk(clk),
                      .reset(reset),
                      .r(and2n_inst2_o0),
                      .s(task_done_pulse),
                      .q(psw_task_done_internal));

  assign task_done_pulse = and2n_inst5_o0 & 1'b1;
  assign and2n_inst2_o0 = sig_clear_task_done & inverter1n_inst7_o0;
  assign inverter1n_inst7_o0 = ~and2n_inst5_o0;

  incdec_counter #(.width(1), .countby(1))  mlinterface_incdec_counter_inst0(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .inc(psw_start_task_init_internal),
                      .dec(psw_start_task_init_internal),
                      .load(1'b0),
                      .i0(1'b0),
                      .o0(psw_livein_frames_in_use_internal));

  sext #(.inwidth(1), .outwidth(4), .signedflag(0))  sext_inst0(
                      .i0(psw_livein_frames_in_use_internal),
                      .o0(sext_inst0_o0[3 : 0]));

  incdec_counter #(.width(1), .countby(1))  mlinterface_incdec_counter_inst1(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .inc(psw_start_task_init_internal),
                      .dec(and2n_inst5_o0),
                      .load(1'b0),
                      .i0(1'b0),
                      .o0(psw_liveout_frames_in_use_internal));

  sext #(.inwidth(1), .outwidth(4), .signedflag(0))  sext_inst1(
                      .i0(psw_liveout_frames_in_use_internal),
                      .o0(sext_inst1_o0[3 : 0]));

  equal #(.width(1))  equal_inst0(
                      .i0(psw_livein_frames_in_use_internal),
                      .i1(1'b0),
                      .o0(equal_inst0_o0));

  equal #(.width(1))  equal_inst1(
                      .i0(psw_liveout_frames_in_use_internal),
                      .i1(1'b0),
                      .o0(equal_inst1_o0));

  assign psw_idle_internal = equal_inst0_o0 & equal_inst1_o0;
  assign psw_released_internal = multiloop_rsflipflop_noinit_inst3_q | psw_start_task_init_internal;
  assign psw_busy_internal = multiloop_rsflipflop_noinit_inst2_q | psw_start_task_init_internal;

  sregn_noinit #(.width(1))  pulsereg_sastatus_0(
                      .clk(clk),
                      .reset(reset),
                      .enable(paw_0_stallbar_out),
                      .i0(inverter1n_inst8_o0),
                      .o0(pulsereg_sastatus_0_o0));

  assign inverter1n_inst8_o0 = ~paw_0_status;
  assign and2n_inst4_o0 = paw_0_status & pulsereg_sastatus_0_o0;

  sregn_noinit #(.width(1))  sregn_noinit_inst5_dly(
                      .clk(clk),
                      .reset(reset),
                      .enable(1'b1),
                      .i0(and2n_inst4_o0),
                      .o0(sregn_noinit_inst5_dly_o0));

  assign psw_sa_0_stalling_internal = ~paw_0_stallbar_out;

  rsflipflop_noinit  multiloop_rsflipflop_noinit_inst2(
                      .clk(clk),
                      .reset(reset),
                      .r(and2n_inst6_o0),
                      .s(psw_start_task_init_internal),
                      .q(multiloop_rsflipflop_noinit_inst2_q));

  rsflipflop_noinit  multiloop_rsflipflop_noinit_inst3(
                      .clk(clk),
                      .reset(reset),
                      .r(and2n_inst7_o0),
                      .s(psw_start_task_init_internal),
                      .q(multiloop_rsflipflop_noinit_inst3_q));

  assign and2n_inst5_o0 = paw_0_status & multiloop_rsflipflop_noinit_inst3_q;
  assign and2n_inst6_o0 = and2n_inst5_o0 & inverter1n_inst10_o0;
  assign inverter1n_inst10_o0 = ~psw_start_task_init_internal;
  assign and2n_inst7_o0 = and2n_inst5_o0 & inverter1n_inst11_o0;
  assign inverter1n_inst11_o0 = ~psw_start_task_init_internal;

  stream_buffer_with_passthru_noreset #(.width(27), .depth(`TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH))  boundary_buf_outstream_dvi_out_dismantle(
                      .clk(clk),
                      .reset(reset),
                      .store_ready(sig_outstream_dvi_out_ready_0),
                      .flush(1'b0),
                      .store_req(boundary_buf_outstream_dvi_out_dismantle_store_req),
                      .load_req(boundary_buf_outstream_dvi_out_dismantle_load_req),
                      .load_ready(paw_0_outstream_dvi_out_req_0),
                      .indata(paw_0_outstream_dvi_out_do_0[26 : 0]),
                      .outdata(boundary_buf_outstream_dvi_out_dismantle_outdata[26 : 0]));


`ifdef TOPLEVEL_test_pattern_generator
// synopsys translate_off
`ifdef CLK_PERIOD
`else
   `define CLK_PERIOD 10.000000
`endif
`ifdef PICO_SYSC_SIM
   `define PICO_PERF_MON
`endif
`ifdef offline_vsim
   `define PICO_PERF_MON
`endif
`ifdef PICO_PERF_MON
   performance_monitor #(.n(1), .m(0),
`ifdef PICO_SYSC_SIM
      .logfilename("online_monitor.log"),
`endif
`ifdef offline_vsim
      .logfilename("transcript_file"),
`endif
      .clk_period(`CLK_PERIOD)
      ) perf_monitor(.clk(clk), .reset(reset), .aborting(1'b0));
`endif // PICO_PERF_MON
// synopsys translate_on


// synopsys translate_off
initial begin
   if (`TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH > 0) begin
`ifdef offline_vsim
      $display("\nWARNING\nWARNING: Output stream 'outstream_dvi_out_dismantle' has a FIFO of depth '%0d'. Note that\n         there could be data inside the FIFO even after the PPA\n         signals task completion.\nEND WARNING\n", `TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH);
`endif // offline_vsim
`ifdef PICO_SYSC_SIM
      $fdisplay(perf_monitor.fileptr, "\nWARNING\nWARNING: Output stream 'outstream_dvi_out_dismantle' has a FIFO of depth '%0d'. Note that\n         there could be data inside the FIFO even after the PPA\n         signals task completion.\nEND WARNING\n", `TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH);
`endif // PICO_SYSC_SIM
   end
end
// synopsys translate_on

// pico offline dump defines:
// synopsys translate_off
`ifdef PICO_DUMP_VCD
      initial begin
                $dumpfile("dump_offline.vcd");
		$dumpvars;
	      end
`endif
`ifdef PICO_DUMP_FSDB
      initial begin
                $fsdbDumpfile("dump_offline.fsdb");
                $fsdbDumpvars ;
              end
`endif
`ifdef PICO_DUMP_VPD
      initial begin
                $vcdplusfile("dump_offline.vpd");
		$vcdpluson;
	      end
`endif
`ifdef PICO_DUMP_TRN
      initial begin
		$recordfile("dump_offline");
		$recordvars;
	      end
`endif
`ifdef PICO_DUMP_VCD_TOP
      initial begin
      		$dumpfile("dump_offline.vcd");
      		$dumpvars (1, test_pattern_generator_testbench.dut.ppa_pico_wrapper_0.ppa_0 );
              end
`endif
`ifdef PICO_DUMP_VCD_PT
      initial begin
      		$dumpfile("dump_offline_pt.vcd");
      		$dumpvars (0, test_pattern_generator_testbench.dut.ppa_pico_wrapper_0.ppa_0 );
              end
`endif
`ifdef PICO_DUMP_VCD_SG
      initial begin
      		$dumpfile("dump_offline_sg.vcd");
      		$dumpvars (0, test_pattern_generator_testbench.dut.ppa_pico_wrapper_0.ppa_0 );
              end
`endif
`ifdef PICO_DUMP_FSDB_PT
      initial begin
                $fsdbDumpfile("dump_offline_pt.fsdb");
                $fsdbDumpvars ;
              end
`endif
`ifdef PICO_DUMP_FSDB_SG
      initial begin
                $fsdbDumpfile("dump_offline_sg.fsdb");
                $fsdbDumpvars ;
              end
`endif
// synopsys translate_on
// pico end offline dump defines:
// 
// pico online dump defines:
// synopsys translate_off
`ifdef PICO_SYSC_SIM
      `ifdef PICO_DUMP_VCD_ONLINE
             initial begin
                       $dumpfile("dump_online.vcd");
		       $dumpvars(0,test_pattern_generator_ppa);
	             end
      `endif
      `ifdef PICO_DUMP_FSDB_ONLINE
             initial begin
                       $fsdbDumpfile("dump_online.fsdb");
                       $fsdbDumpvars (0, test_pattern_generator_ppa );
                     end
      `endif
      `ifdef PICO_DUMP_VPD_ONLINE
             initial begin
                       $vcdplusfile("dump_online.vpd");
		       $vcdpluson;
	             end
      `endif
      `ifdef PICO_DUMP_TRN_ONLINE
             initial begin
		       $recordfile("dump_online");
		       $recordvars(test_pattern_generator_ppa,"depth = 10");
	             end
      `endif
      `ifdef PICO_DUMP_VCD_TOP_ONLINE
       	     initial begin
      		       $dumpfile("dump_online.vcd");
      		       $dumpvars (1, test_pattern_generator_ppa );
                     end
       `endif
      `ifdef PICO_DUMP_VCD_PT_ONLINE
       	     initial begin
      		       $dumpfile("dump_online_pt.vcd");
      		       $dumpvars (0, test_pattern_generator_ppa );
                     end
       `endif
      `ifdef PICO_DUMP_VCD_SG_ONLINE
       	     initial begin
      		       $dumpfile("dump_online_sg.vcd");
      		       $dumpvars (0, test_pattern_generator_ppa );
                     end
       `endif
      `ifdef PICO_DUMP_FSDB_PT_ONLINE
             initial begin
                       $fsdbDumpfile("dump_online_pt.fsdb");
                       $fsdbDumpvars (0, test_pattern_generator_ppa );
                     end
       `endif
      `ifdef PICO_DUMP_FSDB_SG_ONLINE
             initial begin
                       $fsdbDumpfile("dump_online_sg.fsdb");
                       $fsdbDumpvars (0, test_pattern_generator_ppa );
                     end
       `endif
`endif
// synopsys translate_on
// pico end online dump defines
// 
`endif
`ifdef PICO_ASSERTIONS_OFF
`else
 `ifdef ENABLE_ASSERTIONS_IN_RTL
  // pico assertions file instantiation:
  // synopsys translate_off
  test_pattern_generator_ppa_assertions test_pattern_generator_ppa_assertions ();
  // synopsys translate_on
 `endif
`endif
endmodule
// vim: tags=./tags_test_pattern_generator_ppa_v
