/************************************************************************
 *                                                                      *
 * Copyright (c) 2009 Synfora, Inc.  All rights reserved.               *
 *                                                                      *
 * This file contains Confidential Information of Synfora, Inc.         *
 * In addition, certain inventions disclosed in this file may be        *
 * claimed within patents owned or patent applications filed by         *
 * Synfora or third parties.  Any use of Synfora's copyrighted works,   *
 * confidential information, patented inventions, or patent-pending     *
 * inventions is subject to the terms and conditions of your written    *
 * license agreement with Synfora, Inc.                                 *
 * All other use and disclosure is strictly prohibited.                 *
 *                                                                      *
 ************************************************************************/

/* Generated by PICO Extreme FPGA version 09.04 */
/* Target library : xilinx-spartan6-s2 */
/* Target frequency : 100 MHz */

`timescale 1ns / 10 ps

// The following defines named constants used in this file.
`ifdef TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH
`else
`define TEST_PATTERN_GENERATOR_BOUNDARY_BUF_OUTSTREAM_DVI_OUT_DISMANTLE_LENGTH 0
`endif
// End of definitions of named constants

module test_pattern_generator_ppa(
        clk,
        reset,
        start_task_init,
        start_task_final,
        clear_init_done,
        clear_task_done,
        psw_livein_frames_in_use,
        psw_liveout_frames_in_use,
        psw_released,
        psw_sa_0_stalling,
        psw_busy,
        psw_idle,
        psw_init_done,
        psw_task_done,
        rawdatain_hsync_0,
        rawdatain_hblank_0,
        rawdatain_hbporch_0,
        rawdatain_hactive_0,
        rawdatain_vsync_0,
        rawdatain_vblank_0,
        rawdatain_vbporch_0,
        rawdatain_vactive_0,
        rawdatain_hfporch_0,
        rawdatain_vfporch_0,
        outstream_dvi_out_do_0,
        outstream_dvi_out_req_0,
        outstream_dvi_out_ready_0);

  // Module parameters


  // synopsys template

  // Ports

  input  clk;
  input  reset;
  input  start_task_init;
  input  start_task_final;
  input  clear_init_done;
  input  clear_task_done;
  output [3 : 0] psw_livein_frames_in_use;
  output [3 : 0] psw_liveout_frames_in_use;
  output  psw_released;
  output  psw_sa_0_stalling;
  output  psw_busy;
  output  psw_idle;
  output  psw_init_done;
  output  psw_task_done;
  input  rawdatain_hsync_0;
  input [31 : 0] rawdatain_hblank_0;
  input [31 : 0] rawdatain_hbporch_0;
  input [31 : 0] rawdatain_hactive_0;
  input  rawdatain_vsync_0;
  input [31 : 0] rawdatain_vblank_0;
  input [31 : 0] rawdatain_vbporch_0;
  input [31 : 0] rawdatain_vactive_0;
  input [31 : 0] rawdatain_hfporch_0;
  input [31 : 0] rawdatain_vfporch_0;
  output [26 : 0] outstream_dvi_out_do_0;
  output  outstream_dvi_out_req_0;
  input  outstream_dvi_out_ready_0;


endmodule


